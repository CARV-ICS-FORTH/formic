// ===========================================================================
//
//                              FORTH-ICS / CARV
//
//      Licensed under the TAPR Open Hardware License (www.tapr.org/NCL)
//                           Copyright (c) 2010-2012
//
//
// ==========================[ Static Information ]===========================
//
// Author        : Spyros Lyberis
// Abstract      : Full 22-port Crossbar top-level module
//
// =============================[ CVS Variables ]=============================
//
// File name     : $RCSfile: xbar_formic_m8g8.v,v $
// CVS revision  : $Revision: 1.2 $
// Last modified : $Date: 2012/07/03 16:28:58 $
// Last author   : $Author: lyberis $
//
// ===========================================================================

`timescale 1ns/1ps

module xbar_formic_m8g8 (
  
  // Clock and reset
  input         clk_xbar,
  input         rst_xbar,

  // Static configuration
  input   [7:0] i_board_id,

  // Port #00 interface
  output  [2:0] o_port00_out_enq,
  output  [5:0] o_port00_out_offset,
  output        o_port00_out_eop,
  output [15:0] o_port00_out_data,
  input   [2:0] i_port00_out_full,
  input   [2:0] i_port00_out_packets_vc0,
  input   [2:0] i_port00_out_packets_vc1,
  input   [2:0] i_port00_out_packets_vc2,
  output  [2:0] o_port00_in_deq,
  output  [5:0] o_port00_in_offset,
  output        o_port00_in_eop,
  input  [15:0] i_port00_in_data,
  input   [2:0] i_port00_in_empty,

  // Port #01 interface
  output  [2:0] o_port01_out_enq,
  output  [5:0] o_port01_out_offset,
  output        o_port01_out_eop,
  output [15:0] o_port01_out_data,
  input   [2:0] i_port01_out_full,
  input   [2:0] i_port01_out_packets_vc0,
  input   [2:0] i_port01_out_packets_vc1,
  input   [2:0] i_port01_out_packets_vc2,
  output  [2:0] o_port01_in_deq,
  output  [5:0] o_port01_in_offset,
  output        o_port01_in_eop,
  input  [15:0] i_port01_in_data,
  input   [2:0] i_port01_in_empty,

  // Port #02 interface
  output  [2:0] o_port02_out_enq,
  output  [5:0] o_port02_out_offset,
  output        o_port02_out_eop,
  output [15:0] o_port02_out_data,
  input   [2:0] i_port02_out_full,
  input   [2:0] i_port02_out_packets_vc0,
  input   [2:0] i_port02_out_packets_vc1,
  input   [2:0] i_port02_out_packets_vc2,
  output  [2:0] o_port02_in_deq,
  output  [5:0] o_port02_in_offset,
  output        o_port02_in_eop,
  input  [15:0] i_port02_in_data,
  input   [2:0] i_port02_in_empty,

  // Port #03 interface
  output  [2:0] o_port03_out_enq,
  output  [5:0] o_port03_out_offset,
  output        o_port03_out_eop,
  output [15:0] o_port03_out_data,
  input   [2:0] i_port03_out_full,
  input   [2:0] i_port03_out_packets_vc0,
  input   [2:0] i_port03_out_packets_vc1,
  input   [2:0] i_port03_out_packets_vc2,
  output  [2:0] o_port03_in_deq,
  output  [5:0] o_port03_in_offset,
  output        o_port03_in_eop,
  input  [15:0] i_port03_in_data,
  input   [2:0] i_port03_in_empty,

  // Port #04 interface
  output  [2:0] o_port04_out_enq,
  output  [5:0] o_port04_out_offset,
  output        o_port04_out_eop,
  output [15:0] o_port04_out_data,
  input   [2:0] i_port04_out_full,
  input   [2:0] i_port04_out_packets_vc0,
  input   [2:0] i_port04_out_packets_vc1,
  input   [2:0] i_port04_out_packets_vc2,
  output  [2:0] o_port04_in_deq,
  output  [5:0] o_port04_in_offset,
  output        o_port04_in_eop,
  input  [15:0] i_port04_in_data,
  input   [2:0] i_port04_in_empty,

  // Port #05 interface
  output  [2:0] o_port05_out_enq,
  output  [5:0] o_port05_out_offset,
  output        o_port05_out_eop,
  output [15:0] o_port05_out_data,
  input   [2:0] i_port05_out_full,
  input   [2:0] i_port05_out_packets_vc0,
  input   [2:0] i_port05_out_packets_vc1,
  input   [2:0] i_port05_out_packets_vc2,
  output  [2:0] o_port05_in_deq,
  output  [5:0] o_port05_in_offset,
  output        o_port05_in_eop,
  input  [15:0] i_port05_in_data,
  input   [2:0] i_port05_in_empty,

  // Port #06 interface
  output  [2:0] o_port06_out_enq,
  output  [5:0] o_port06_out_offset,
  output        o_port06_out_eop,
  output [15:0] o_port06_out_data,
  input   [2:0] i_port06_out_full,
  input   [2:0] i_port06_out_packets_vc0,
  input   [2:0] i_port06_out_packets_vc1,
  input   [2:0] i_port06_out_packets_vc2,
  output  [2:0] o_port06_in_deq,
  output  [5:0] o_port06_in_offset,
  output        o_port06_in_eop,
  input  [15:0] i_port06_in_data,
  input   [2:0] i_port06_in_empty,

  // Port #07 interface
  output  [2:0] o_port07_out_enq,
  output  [5:0] o_port07_out_offset,
  output        o_port07_out_eop,
  output [15:0] o_port07_out_data,
  input   [2:0] i_port07_out_full,
  input   [2:0] i_port07_out_packets_vc0,
  input   [2:0] i_port07_out_packets_vc1,
  input   [2:0] i_port07_out_packets_vc2,
  output  [2:0] o_port07_in_deq,
  output  [5:0] o_port07_in_offset,
  output        o_port07_in_eop,
  input  [15:0] i_port07_in_data,
  input   [2:0] i_port07_in_empty,

  // Port #08 interface
  output  [2:0] o_port08_out_enq,
  output  [5:0] o_port08_out_offset,
  output        o_port08_out_eop,
  output [15:0] o_port08_out_data,
  input   [2:0] i_port08_out_full,
  input   [2:0] i_port08_out_packets_vc0,
  input   [2:0] i_port08_out_packets_vc1,
  input   [2:0] i_port08_out_packets_vc2,
  output  [2:0] o_port08_in_deq,
  output  [5:0] o_port08_in_offset,
  output        o_port08_in_eop,
  input  [15:0] i_port08_in_data,
  input   [2:0] i_port08_in_empty,

  // Port #09 interface
  output  [2:0] o_port09_out_enq,
  output  [5:0] o_port09_out_offset,
  output        o_port09_out_eop,
  output [15:0] o_port09_out_data,
  input   [2:0] i_port09_out_full,
  input   [2:0] i_port09_out_packets_vc0,
  input   [2:0] i_port09_out_packets_vc1,
  input   [2:0] i_port09_out_packets_vc2,
  output  [2:0] o_port09_in_deq,
  output  [5:0] o_port09_in_offset,
  output        o_port09_in_eop,
  input  [15:0] i_port09_in_data,
  input   [2:0] i_port09_in_empty,

  // Port #10 interface
  output  [2:0] o_port10_out_enq,
  output  [5:0] o_port10_out_offset,
  output        o_port10_out_eop,
  output [15:0] o_port10_out_data,
  input   [2:0] i_port10_out_full,
  input   [2:0] i_port10_out_packets_vc0,
  input   [2:0] i_port10_out_packets_vc1,
  input   [2:0] i_port10_out_packets_vc2,
  output  [2:0] o_port10_in_deq,
  output  [5:0] o_port10_in_offset,
  output        o_port10_in_eop,
  input  [15:0] i_port10_in_data,
  input   [2:0] i_port10_in_empty,

  // Port #11 interface
  output  [2:0] o_port11_out_enq,
  output  [5:0] o_port11_out_offset,
  output        o_port11_out_eop,
  output [15:0] o_port11_out_data,
  input   [2:0] i_port11_out_full,
  input   [2:0] i_port11_out_packets_vc0,
  input   [2:0] i_port11_out_packets_vc1,
  input   [2:0] i_port11_out_packets_vc2,
  output  [2:0] o_port11_in_deq,
  output  [5:0] o_port11_in_offset,
  output        o_port11_in_eop,
  input  [15:0] i_port11_in_data,
  input   [2:0] i_port11_in_empty,

  // Port #12 interface
  output  [2:0] o_port12_out_enq,
  output  [5:0] o_port12_out_offset,
  output        o_port12_out_eop,
  output [15:0] o_port12_out_data,
  input   [2:0] i_port12_out_full,
  input   [2:0] i_port12_out_packets_vc0,
  input   [2:0] i_port12_out_packets_vc1,
  input   [2:0] i_port12_out_packets_vc2,
  output  [2:0] o_port12_in_deq,
  output  [5:0] o_port12_in_offset,
  output        o_port12_in_eop,
  input  [15:0] i_port12_in_data,
  input   [2:0] i_port12_in_empty,

  // Port #13 interface
  output  [2:0] o_port13_out_enq,
  output  [5:0] o_port13_out_offset,
  output        o_port13_out_eop,
  output [15:0] o_port13_out_data,
  input   [2:0] i_port13_out_full,
  input   [2:0] i_port13_out_packets_vc0,
  input   [2:0] i_port13_out_packets_vc1,
  input   [2:0] i_port13_out_packets_vc2,
  output  [2:0] o_port13_in_deq,
  output  [5:0] o_port13_in_offset,
  output        o_port13_in_eop,
  input  [15:0] i_port13_in_data,
  input   [2:0] i_port13_in_empty,

  // Port #14 interface
  output  [2:0] o_port14_out_enq,
  output  [5:0] o_port14_out_offset,
  output        o_port14_out_eop,
  output [15:0] o_port14_out_data,
  input   [2:0] i_port14_out_full,
  input   [2:0] i_port14_out_packets_vc0,
  input   [2:0] i_port14_out_packets_vc1,
  input   [2:0] i_port14_out_packets_vc2,
  output  [2:0] o_port14_in_deq,
  output  [5:0] o_port14_in_offset,
  output        o_port14_in_eop,
  input  [15:0] i_port14_in_data,
  input   [2:0] i_port14_in_empty,

  // Port #15 interface
  output  [2:0] o_port15_out_enq,
  output  [5:0] o_port15_out_offset,
  output        o_port15_out_eop,
  output [15:0] o_port15_out_data,
  input   [2:0] i_port15_out_full,
  input   [2:0] i_port15_out_packets_vc0,
  input   [2:0] i_port15_out_packets_vc1,
  input   [2:0] i_port15_out_packets_vc2,
  output  [2:0] o_port15_in_deq,
  output  [5:0] o_port15_in_offset,
  output        o_port15_in_eop,
  input  [15:0] i_port15_in_data,
  input   [2:0] i_port15_in_empty,

  // Port #16 interface
  output  [2:0] o_port16_out_enq,
  output  [5:0] o_port16_out_offset,
  output        o_port16_out_eop,
  output [15:0] o_port16_out_data,
  input   [2:0] i_port16_out_full,
  input   [2:0] i_port16_out_packets_vc0,
  input   [2:0] i_port16_out_packets_vc1,
  input   [2:0] i_port16_out_packets_vc2,
  output  [2:0] o_port16_in_deq,
  output  [5:0] o_port16_in_offset,
  output        o_port16_in_eop,
  input  [15:0] i_port16_in_data,
  input   [2:0] i_port16_in_empty,

  // Port #17 interface
  output  [2:0] o_port17_out_enq,
  output  [5:0] o_port17_out_offset,
  output        o_port17_out_eop,
  output [15:0] o_port17_out_data,
  input   [2:0] i_port17_out_full,
  input   [2:0] i_port17_out_packets_vc0,
  input   [2:0] i_port17_out_packets_vc1,
  input   [2:0] i_port17_out_packets_vc2,
  output  [2:0] o_port17_in_deq,
  output  [5:0] o_port17_in_offset,
  output        o_port17_in_eop,
  input  [15:0] i_port17_in_data,
  input   [2:0] i_port17_in_empty,

  // Port #18 interface
  output  [2:0] o_port18_out_enq,
  output  [5:0] o_port18_out_offset,
  output        o_port18_out_eop,
  output [15:0] o_port18_out_data,
  input   [2:0] i_port18_out_full,
  input   [2:0] i_port18_out_packets_vc0,
  input   [2:0] i_port18_out_packets_vc1,
  input   [2:0] i_port18_out_packets_vc2,
  output  [2:0] o_port18_in_deq,
  output  [5:0] o_port18_in_offset,
  output        o_port18_in_eop,
  input  [15:0] i_port18_in_data,
  input   [2:0] i_port18_in_empty,

  // Port #19 interface
  output  [2:0] o_port19_out_enq,
  output  [5:0] o_port19_out_offset,
  output        o_port19_out_eop,
  output [15:0] o_port19_out_data,
  input   [2:0] i_port19_out_full,
  input   [2:0] i_port19_out_packets_vc0,
  input   [2:0] i_port19_out_packets_vc1,
  input   [2:0] i_port19_out_packets_vc2,
  output  [2:0] o_port19_in_deq,
  output  [5:0] o_port19_in_offset,
  output        o_port19_in_eop,
  input  [15:0] i_port19_in_data,
  input   [2:0] i_port19_in_empty,

  // Port #20 interface
  output  [2:0] o_port20_out_enq,
  output  [5:0] o_port20_out_offset,
  output        o_port20_out_eop,
  output [15:0] o_port20_out_data,
  input   [2:0] i_port20_out_full,
  input   [2:0] i_port20_out_packets_vc0,
  input   [2:0] i_port20_out_packets_vc1,
  input   [2:0] i_port20_out_packets_vc2,
  output  [2:0] o_port20_in_deq,
  output  [5:0] o_port20_in_offset,
  output        o_port20_in_eop,
  input  [15:0] i_port20_in_data,
  input   [2:0] i_port20_in_empty,

  // Port #21 interface
  output  [2:0] o_port21_out_enq,
  output  [5:0] o_port21_out_offset,
  output        o_port21_out_eop,
  output [15:0] o_port21_out_data,
  input   [2:0] i_port21_out_full,
  input   [2:0] i_port21_out_packets_vc0,
  input   [2:0] i_port21_out_packets_vc1,
  input   [2:0] i_port21_out_packets_vc2,
  output  [2:0] o_port21_in_deq,
  output  [5:0] o_port21_in_offset,
  output        o_port21_in_eop,
  input  [15:0] i_port21_in_data,
  input   [2:0] i_port21_in_empty
);

  // ==========================================================================
  // Wires
  // ==========================================================================
  wire [21:0] arbin00_req0;
  wire [21:0] arbin00_req1;
  wire [21:0] arbin00_req2;
  wire [21:0] arbin00_gnt0;
  wire [21:0] arbin00_gnt1;
  wire [21:0] arbin00_gnt2;
  wire [15:0] arbin00_data;

  wire [21:0] arbin01_req0;
  wire [21:0] arbin01_req1;
  wire [21:0] arbin01_req2;
  wire [21:0] arbin01_gnt0;
  wire [21:0] arbin01_gnt1;
  wire [21:0] arbin01_gnt2;
  wire [15:0] arbin01_data;

  wire [21:0] arbin02_req0;
  wire [21:0] arbin02_req1;
  wire [21:0] arbin02_req2;
  wire [21:0] arbin02_gnt0;
  wire [21:0] arbin02_gnt1;
  wire [21:0] arbin02_gnt2;
  wire [15:0] arbin02_data;

  wire [21:0] arbin03_req0;
  wire [21:0] arbin03_req1;
  wire [21:0] arbin03_req2;
  wire [21:0] arbin03_gnt0;
  wire [21:0] arbin03_gnt1;
  wire [21:0] arbin03_gnt2;
  wire [15:0] arbin03_data;

  wire [21:0] arbin04_req0;
  wire [21:0] arbin04_req1;
  wire [21:0] arbin04_req2;
  wire [21:0] arbin04_gnt0;
  wire [21:0] arbin04_gnt1;
  wire [21:0] arbin04_gnt2;
  wire [15:0] arbin04_data;

  wire [21:0] arbin05_req0;
  wire [21:0] arbin05_req1;
  wire [21:0] arbin05_req2;
  wire [21:0] arbin05_gnt0;
  wire [21:0] arbin05_gnt1;
  wire [21:0] arbin05_gnt2;
  wire [15:0] arbin05_data;

  wire [21:0] arbin06_req0;
  wire [21:0] arbin06_req1;
  wire [21:0] arbin06_req2;
  wire [21:0] arbin06_gnt0;
  wire [21:0] arbin06_gnt1;
  wire [21:0] arbin06_gnt2;
  wire [15:0] arbin06_data;

  wire [21:0] arbin07_req0;
  wire [21:0] arbin07_req1;
  wire [21:0] arbin07_req2;
  wire [21:0] arbin07_gnt0;
  wire [21:0] arbin07_gnt1;
  wire [21:0] arbin07_gnt2;
  wire [15:0] arbin07_data;

  wire [21:0] arbin08_req0;
  wire [21:0] arbin08_req1;
  wire [21:0] arbin08_req2;
  wire [21:0] arbin08_gnt0;
  wire [21:0] arbin08_gnt1;
  wire [21:0] arbin08_gnt2;
  wire [15:0] arbin08_data;

  wire [21:0] arbin09_req0;
  wire [21:0] arbin09_req1;
  wire [21:0] arbin09_req2;
  wire [21:0] arbin09_gnt0;
  wire [21:0] arbin09_gnt1;
  wire [21:0] arbin09_gnt2;
  wire [15:0] arbin09_data;

  wire [21:0] arbin10_req0;
  wire [21:0] arbin10_req1;
  wire [21:0] arbin10_req2;
  wire [21:0] arbin10_gnt0;
  wire [21:0] arbin10_gnt1;
  wire [21:0] arbin10_gnt2;
  wire [15:0] arbin10_data;

  wire [21:0] arbin11_req0;
  wire [21:0] arbin11_req1;
  wire [21:0] arbin11_req2;
  wire [21:0] arbin11_gnt0;
  wire [21:0] arbin11_gnt1;
  wire [21:0] arbin11_gnt2;
  wire [15:0] arbin11_data;

  wire [21:0] arbin12_req0;
  wire [21:0] arbin12_req1;
  wire [21:0] arbin12_req2;
  wire [21:0] arbin12_gnt0;
  wire [21:0] arbin12_gnt1;
  wire [21:0] arbin12_gnt2;
  wire [15:0] arbin12_data;

  wire [21:0] arbin13_req0;
  wire [21:0] arbin13_req1;
  wire [21:0] arbin13_req2;
  wire [21:0] arbin13_gnt0;
  wire [21:0] arbin13_gnt1;
  wire [21:0] arbin13_gnt2;
  wire [15:0] arbin13_data;

  wire [21:0] arbin14_req0;
  wire [21:0] arbin14_req1;
  wire [21:0] arbin14_req2;
  wire [21:0] arbin14_gnt0;
  wire [21:0] arbin14_gnt1;
  wire [21:0] arbin14_gnt2;
  wire [15:0] arbin14_data;

  wire [21:0] arbin15_req0;
  wire [21:0] arbin15_req1;
  wire [21:0] arbin15_req2;
  wire [21:0] arbin15_gnt0;
  wire [21:0] arbin15_gnt1;
  wire [21:0] arbin15_gnt2;
  wire [15:0] arbin15_data;

  wire [21:0] arbin16_req0;
  wire [21:0] arbin16_req1;
  wire [21:0] arbin16_req2;
  wire [21:0] arbin16_gnt0;
  wire [21:0] arbin16_gnt1;
  wire [21:0] arbin16_gnt2;
  wire [15:0] arbin16_data;

  wire [21:0] arbin17_req0;
  wire [21:0] arbin17_req1;
  wire [21:0] arbin17_req2;
  wire [21:0] arbin17_gnt0;
  wire [21:0] arbin17_gnt1;
  wire [21:0] arbin17_gnt2;
  wire [15:0] arbin17_data;

  wire [21:0] arbin18_req0;
  wire [21:0] arbin18_req1;
  wire [21:0] arbin18_req2;
  wire [21:0] arbin18_gnt0;
  wire [21:0] arbin18_gnt1;
  wire [21:0] arbin18_gnt2;
  wire [15:0] arbin18_data;

  wire [21:0] arbin19_req0;
  wire [21:0] arbin19_req1;
  wire [21:0] arbin19_req2;
  wire [21:0] arbin19_gnt0;
  wire [21:0] arbin19_gnt1;
  wire [21:0] arbin19_gnt2;
  wire [15:0] arbin19_data;

  wire [21:0] arbin20_req0;
  wire [21:0] arbin20_req1;
  wire [21:0] arbin20_req2;
  wire [21:0] arbin20_gnt0;
  wire [21:0] arbin20_gnt1;
  wire [21:0] arbin20_gnt2;
  wire [15:0] arbin20_data;

  wire [21:0] arbin21_req0;
  wire [21:0] arbin21_req1;
  wire [21:0] arbin21_req2;
  wire [21:0] arbin21_gnt0;
  wire [21:0] arbin21_gnt1;
  wire [21:0] arbin21_gnt2;
  wire [15:0] arbin21_data;


  wire [21:0] arbout00_req0;
  wire [21:0] arbout00_req1;
  wire [21:0] arbout00_req2;
  wire [21:0] arbout00_gnt0;
  wire [21:0] arbout00_gnt1;
  wire [21:0] arbout00_gnt2;
  wire  [4:0] arbout00_mux_sel;
  wire [15:0] arbout00_data;

  wire [21:0] arbout01_req0;
  wire [21:0] arbout01_req1;
  wire [21:0] arbout01_req2;
  wire [21:0] arbout01_gnt0;
  wire [21:0] arbout01_gnt1;
  wire [21:0] arbout01_gnt2;
  wire  [4:0] arbout01_mux_sel;
  wire [15:0] arbout01_data;

  wire [21:0] arbout02_req0;
  wire [21:0] arbout02_req1;
  wire [21:0] arbout02_req2;
  wire [21:0] arbout02_gnt0;
  wire [21:0] arbout02_gnt1;
  wire [21:0] arbout02_gnt2;
  wire  [4:0] arbout02_mux_sel;
  wire [15:0] arbout02_data;

  wire [21:0] arbout03_req0;
  wire [21:0] arbout03_req1;
  wire [21:0] arbout03_req2;
  wire [21:0] arbout03_gnt0;
  wire [21:0] arbout03_gnt1;
  wire [21:0] arbout03_gnt2;
  wire  [4:0] arbout03_mux_sel;
  wire [15:0] arbout03_data;

  wire [21:0] arbout04_req0;
  wire [21:0] arbout04_req1;
  wire [21:0] arbout04_req2;
  wire [21:0] arbout04_gnt0;
  wire [21:0] arbout04_gnt1;
  wire [21:0] arbout04_gnt2;
  wire  [4:0] arbout04_mux_sel;
  wire [15:0] arbout04_data;

  wire [21:0] arbout05_req0;
  wire [21:0] arbout05_req1;
  wire [21:0] arbout05_req2;
  wire [21:0] arbout05_gnt0;
  wire [21:0] arbout05_gnt1;
  wire [21:0] arbout05_gnt2;
  wire  [4:0] arbout05_mux_sel;
  wire [15:0] arbout05_data;

  wire [21:0] arbout06_req0;
  wire [21:0] arbout06_req1;
  wire [21:0] arbout06_req2;
  wire [21:0] arbout06_gnt0;
  wire [21:0] arbout06_gnt1;
  wire [21:0] arbout06_gnt2;
  wire  [4:0] arbout06_mux_sel;
  wire [15:0] arbout06_data;

  wire [21:0] arbout07_req0;
  wire [21:0] arbout07_req1;
  wire [21:0] arbout07_req2;
  wire [21:0] arbout07_gnt0;
  wire [21:0] arbout07_gnt1;
  wire [21:0] arbout07_gnt2;
  wire  [4:0] arbout07_mux_sel;
  wire [15:0] arbout07_data;

  wire [21:0] arbout08_req0;
  wire [21:0] arbout08_req1;
  wire [21:0] arbout08_req2;
  wire [21:0] arbout08_gnt0;
  wire [21:0] arbout08_gnt1;
  wire [21:0] arbout08_gnt2;
  wire  [4:0] arbout08_mux_sel;
  wire [15:0] arbout08_data;

  wire [21:0] arbout09_req0;
  wire [21:0] arbout09_req1;
  wire [21:0] arbout09_req2;
  wire [21:0] arbout09_gnt0;
  wire [21:0] arbout09_gnt1;
  wire [21:0] arbout09_gnt2;
  wire  [4:0] arbout09_mux_sel;
  wire [15:0] arbout09_data;

  wire [21:0] arbout10_req0;
  wire [21:0] arbout10_req1;
  wire [21:0] arbout10_req2;
  wire [21:0] arbout10_gnt0;
  wire [21:0] arbout10_gnt1;
  wire [21:0] arbout10_gnt2;
  wire  [4:0] arbout10_mux_sel;
  wire [15:0] arbout10_data;

  wire [21:0] arbout11_req0;
  wire [21:0] arbout11_req1;
  wire [21:0] arbout11_req2;
  wire [21:0] arbout11_gnt0;
  wire [21:0] arbout11_gnt1;
  wire [21:0] arbout11_gnt2;
  wire  [4:0] arbout11_mux_sel;
  wire [15:0] arbout11_data;

  wire [21:0] arbout12_req0;
  wire [21:0] arbout12_req1;
  wire [21:0] arbout12_req2;
  wire [21:0] arbout12_gnt0;
  wire [21:0] arbout12_gnt1;
  wire [21:0] arbout12_gnt2;
  wire  [4:0] arbout12_mux_sel;
  wire [15:0] arbout12_data;

  wire [21:0] arbout13_req0;
  wire [21:0] arbout13_req1;
  wire [21:0] arbout13_req2;
  wire [21:0] arbout13_gnt0;
  wire [21:0] arbout13_gnt1;
  wire [21:0] arbout13_gnt2;
  wire  [4:0] arbout13_mux_sel;
  wire [15:0] arbout13_data;

  wire [21:0] arbout14_req0;
  wire [21:0] arbout14_req1;
  wire [21:0] arbout14_req2;
  wire [21:0] arbout14_gnt0;
  wire [21:0] arbout14_gnt1;
  wire [21:0] arbout14_gnt2;
  wire  [4:0] arbout14_mux_sel;
  wire [15:0] arbout14_data;

  wire [21:0] arbout15_req0;
  wire [21:0] arbout15_req1;
  wire [21:0] arbout15_req2;
  wire [21:0] arbout15_gnt0;
  wire [21:0] arbout15_gnt1;
  wire [21:0] arbout15_gnt2;
  wire  [4:0] arbout15_mux_sel;
  wire [15:0] arbout15_data;

  wire [21:0] arbout16_req0;
  wire [21:0] arbout16_req1;
  wire [21:0] arbout16_req2;
  wire [21:0] arbout16_gnt0;
  wire [21:0] arbout16_gnt1;
  wire [21:0] arbout16_gnt2;
  wire  [4:0] arbout16_mux_sel;
  wire [15:0] arbout16_data;

  wire [21:0] arbout17_req0;
  wire [21:0] arbout17_req1;
  wire [21:0] arbout17_req2;
  wire [21:0] arbout17_gnt0;
  wire [21:0] arbout17_gnt1;
  wire [21:0] arbout17_gnt2;
  wire  [4:0] arbout17_mux_sel;
  wire [15:0] arbout17_data;

  wire [21:0] arbout18_req0;
  wire [21:0] arbout18_req1;
  wire [21:0] arbout18_req2;
  wire [21:0] arbout18_gnt0;
  wire [21:0] arbout18_gnt1;
  wire [21:0] arbout18_gnt2;
  wire  [4:0] arbout18_mux_sel;
  wire [15:0] arbout18_data;

  wire [21:0] arbout19_req0;
  wire [21:0] arbout19_req1;
  wire [21:0] arbout19_req2;
  wire [21:0] arbout19_gnt0;
  wire [21:0] arbout19_gnt1;
  wire [21:0] arbout19_gnt2;
  wire  [4:0] arbout19_mux_sel;
  wire [15:0] arbout19_data;

  wire [21:0] arbout20_req0;
  wire [21:0] arbout20_req1;
  wire [21:0] arbout20_req2;
  wire [21:0] arbout20_gnt0;
  wire [21:0] arbout20_gnt1;
  wire [21:0] arbout20_gnt2;
  wire  [4:0] arbout20_mux_sel;
  wire [15:0] arbout20_data;

  wire [21:0] arbout21_req0;
  wire [21:0] arbout21_req1;
  wire [21:0] arbout21_req2;
  wire [21:0] arbout21_gnt0;
  wire [21:0] arbout21_gnt1;
  wire [21:0] arbout21_gnt2;
  wire  [4:0] arbout21_mux_sel;
  wire [15:0] arbout21_data;


  // ==========================================================================
  // Input Arbiters
  // ==========================================================================
  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i00_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port00_in_deq ), 
    .o_fifo_offset          ( o_port00_in_offset ),
    .o_fifo_eop             ( o_port00_in_eop ), 
    .i_fifo_data            ( i_port00_in_data ),
    .i_fifo_empty           ( i_port00_in_empty ),
    .o_req0                 ( arbin00_req0 ),
    .o_req1                 ( arbin00_req1 ),
    .o_req2                 ( arbin00_req2 ),
    .i_gnt0                 ( arbin00_gnt0 ),
    .i_gnt1                 ( arbin00_gnt1 ),
    .i_gnt2                 ( arbin00_gnt2 ),
    .o_data                 ( arbin00_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i01_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port01_in_deq ), 
    .o_fifo_offset          ( o_port01_in_offset ),
    .o_fifo_eop             ( o_port01_in_eop ), 
    .i_fifo_data            ( i_port01_in_data ),
    .i_fifo_empty           ( i_port01_in_empty ),
    .o_req0                 ( arbin01_req0 ),
    .o_req1                 ( arbin01_req1 ),
    .o_req2                 ( arbin01_req2 ),
    .i_gnt0                 ( arbin01_gnt0 ),
    .i_gnt1                 ( arbin01_gnt1 ),
    .i_gnt2                 ( arbin01_gnt2 ),
    .o_data                 ( arbin01_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i02_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port02_in_deq ), 
    .o_fifo_offset          ( o_port02_in_offset ),
    .o_fifo_eop             ( o_port02_in_eop ), 
    .i_fifo_data            ( i_port02_in_data ),
    .i_fifo_empty           ( i_port02_in_empty ),
    .o_req0                 ( arbin02_req0 ),
    .o_req1                 ( arbin02_req1 ),
    .o_req2                 ( arbin02_req2 ),
    .i_gnt0                 ( arbin02_gnt0 ),
    .i_gnt1                 ( arbin02_gnt1 ),
    .i_gnt2                 ( arbin02_gnt2 ),
    .o_data                 ( arbin02_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i03_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port03_in_deq ), 
    .o_fifo_offset          ( o_port03_in_offset ),
    .o_fifo_eop             ( o_port03_in_eop ), 
    .i_fifo_data            ( i_port03_in_data ),
    .i_fifo_empty           ( i_port03_in_empty ),
    .o_req0                 ( arbin03_req0 ),
    .o_req1                 ( arbin03_req1 ),
    .o_req2                 ( arbin03_req2 ),
    .i_gnt0                 ( arbin03_gnt0 ),
    .i_gnt1                 ( arbin03_gnt1 ),
    .i_gnt2                 ( arbin03_gnt2 ),
    .o_data                 ( arbin03_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i04_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port04_in_deq ), 
    .o_fifo_offset          ( o_port04_in_offset ),
    .o_fifo_eop             ( o_port04_in_eop ), 
    .i_fifo_data            ( i_port04_in_data ),
    .i_fifo_empty           ( i_port04_in_empty ),
    .o_req0                 ( arbin04_req0 ),
    .o_req1                 ( arbin04_req1 ),
    .o_req2                 ( arbin04_req2 ),
    .i_gnt0                 ( arbin04_gnt0 ),
    .i_gnt1                 ( arbin04_gnt1 ),
    .i_gnt2                 ( arbin04_gnt2 ),
    .o_data                 ( arbin04_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i05_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port05_in_deq ), 
    .o_fifo_offset          ( o_port05_in_offset ),
    .o_fifo_eop             ( o_port05_in_eop ), 
    .i_fifo_data            ( i_port05_in_data ),
    .i_fifo_empty           ( i_port05_in_empty ),
    .o_req0                 ( arbin05_req0 ),
    .o_req1                 ( arbin05_req1 ),
    .o_req2                 ( arbin05_req2 ),
    .i_gnt0                 ( arbin05_gnt0 ),
    .i_gnt1                 ( arbin05_gnt1 ),
    .i_gnt2                 ( arbin05_gnt2 ),
    .o_data                 ( arbin05_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i06_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port06_in_deq ), 
    .o_fifo_offset          ( o_port06_in_offset ),
    .o_fifo_eop             ( o_port06_in_eop ), 
    .i_fifo_data            ( i_port06_in_data ),
    .i_fifo_empty           ( i_port06_in_empty ),
    .o_req0                 ( arbin06_req0 ),
    .o_req1                 ( arbin06_req1 ),
    .o_req2                 ( arbin06_req2 ),
    .i_gnt0                 ( arbin06_gnt0 ),
    .i_gnt1                 ( arbin06_gnt1 ),
    .i_gnt2                 ( arbin06_gnt2 ),
    .o_data                 ( arbin06_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i07_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port07_in_deq ), 
    .o_fifo_offset          ( o_port07_in_offset ),
    .o_fifo_eop             ( o_port07_in_eop ), 
    .i_fifo_data            ( i_port07_in_data ),
    .i_fifo_empty           ( i_port07_in_empty ),
    .o_req0                 ( arbin07_req0 ),
    .o_req1                 ( arbin07_req1 ),
    .o_req2                 ( arbin07_req2 ),
    .i_gnt0                 ( arbin07_gnt0 ),
    .i_gnt1                 ( arbin07_gnt1 ),
    .i_gnt2                 ( arbin07_gnt2 ),
    .o_data                 ( arbin07_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i08_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port08_in_deq ), 
    .o_fifo_offset          ( o_port08_in_offset ),
    .o_fifo_eop             ( o_port08_in_eop ), 
    .i_fifo_data            ( i_port08_in_data ),
    .i_fifo_empty           ( i_port08_in_empty ),
    .o_req0                 ( arbin08_req0 ),
    .o_req1                 ( arbin08_req1 ),
    .o_req2                 ( arbin08_req2 ),
    .i_gnt0                 ( arbin08_gnt0 ),
    .i_gnt1                 ( arbin08_gnt1 ),
    .i_gnt2                 ( arbin08_gnt2 ),
    .o_data                 ( arbin08_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i09_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port09_in_deq ), 
    .o_fifo_offset          ( o_port09_in_offset ),
    .o_fifo_eop             ( o_port09_in_eop ), 
    .i_fifo_data            ( i_port09_in_data ),
    .i_fifo_empty           ( i_port09_in_empty ),
    .o_req0                 ( arbin09_req0 ),
    .o_req1                 ( arbin09_req1 ),
    .o_req2                 ( arbin09_req2 ),
    .i_gnt0                 ( arbin09_gnt0 ),
    .i_gnt1                 ( arbin09_gnt1 ),
    .i_gnt2                 ( arbin09_gnt2 ),
    .o_data                 ( arbin09_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i10_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port10_in_deq ), 
    .o_fifo_offset          ( o_port10_in_offset ),
    .o_fifo_eop             ( o_port10_in_eop ), 
    .i_fifo_data            ( i_port10_in_data ),
    .i_fifo_empty           ( i_port10_in_empty ),
    .o_req0                 ( arbin10_req0 ),
    .o_req1                 ( arbin10_req1 ),
    .o_req2                 ( arbin10_req2 ),
    .i_gnt0                 ( arbin10_gnt0 ),
    .i_gnt1                 ( arbin10_gnt1 ),
    .i_gnt2                 ( arbin10_gnt2 ),
    .o_data                 ( arbin10_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i11_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port11_in_deq ), 
    .o_fifo_offset          ( o_port11_in_offset ),
    .o_fifo_eop             ( o_port11_in_eop ), 
    .i_fifo_data            ( i_port11_in_data ),
    .i_fifo_empty           ( i_port11_in_empty ),
    .o_req0                 ( arbin11_req0 ),
    .o_req1                 ( arbin11_req1 ),
    .o_req2                 ( arbin11_req2 ),
    .i_gnt0                 ( arbin11_gnt0 ),
    .i_gnt1                 ( arbin11_gnt1 ),
    .i_gnt2                 ( arbin11_gnt2 ),
    .o_data                 ( arbin11_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i12_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port12_in_deq ), 
    .o_fifo_offset          ( o_port12_in_offset ),
    .o_fifo_eop             ( o_port12_in_eop ), 
    .i_fifo_data            ( i_port12_in_data ),
    .i_fifo_empty           ( i_port12_in_empty ),
    .o_req0                 ( arbin12_req0 ),
    .o_req1                 ( arbin12_req1 ),
    .o_req2                 ( arbin12_req2 ),
    .i_gnt0                 ( arbin12_gnt0 ),
    .i_gnt1                 ( arbin12_gnt1 ),
    .i_gnt2                 ( arbin12_gnt2 ),
    .o_data                 ( arbin12_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i13_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port13_in_deq ), 
    .o_fifo_offset          ( o_port13_in_offset ),
    .o_fifo_eop             ( o_port13_in_eop ), 
    .i_fifo_data            ( i_port13_in_data ),
    .i_fifo_empty           ( i_port13_in_empty ),
    .o_req0                 ( arbin13_req0 ),
    .o_req1                 ( arbin13_req1 ),
    .o_req2                 ( arbin13_req2 ),
    .i_gnt0                 ( arbin13_gnt0 ),
    .i_gnt1                 ( arbin13_gnt1 ),
    .i_gnt2                 ( arbin13_gnt2 ),
    .o_data                 ( arbin13_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i14_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port14_in_deq ), 
    .o_fifo_offset          ( o_port14_in_offset ),
    .o_fifo_eop             ( o_port14_in_eop ), 
    .i_fifo_data            ( i_port14_in_data ),
    .i_fifo_empty           ( i_port14_in_empty ),
    .o_req0                 ( arbin14_req0 ),
    .o_req1                 ( arbin14_req1 ),
    .o_req2                 ( arbin14_req2 ),
    .i_gnt0                 ( arbin14_gnt0 ),
    .i_gnt1                 ( arbin14_gnt1 ),
    .i_gnt2                 ( arbin14_gnt2 ),
    .o_data                 ( arbin14_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i15_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port15_in_deq ), 
    .o_fifo_offset          ( o_port15_in_offset ),
    .o_fifo_eop             ( o_port15_in_eop ), 
    .i_fifo_data            ( i_port15_in_data ),
    .i_fifo_empty           ( i_port15_in_empty ),
    .o_req0                 ( arbin15_req0 ),
    .o_req1                 ( arbin15_req1 ),
    .o_req2                 ( arbin15_req2 ),
    .i_gnt0                 ( arbin15_gnt0 ),
    .i_gnt1                 ( arbin15_gnt1 ),
    .i_gnt2                 ( arbin15_gnt2 ),
    .o_data                 ( arbin15_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i16_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port16_in_deq ), 
    .o_fifo_offset          ( o_port16_in_offset ),
    .o_fifo_eop             ( o_port16_in_eop ), 
    .i_fifo_data            ( i_port16_in_data ),
    .i_fifo_empty           ( i_port16_in_empty ),
    .o_req0                 ( arbin16_req0 ),
    .o_req1                 ( arbin16_req1 ),
    .o_req2                 ( arbin16_req2 ),
    .i_gnt0                 ( arbin16_gnt0 ),
    .i_gnt1                 ( arbin16_gnt1 ),
    .i_gnt2                 ( arbin16_gnt2 ),
    .o_data                 ( arbin16_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i17_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port17_in_deq ), 
    .o_fifo_offset          ( o_port17_in_offset ),
    .o_fifo_eop             ( o_port17_in_eop ), 
    .i_fifo_data            ( i_port17_in_data ),
    .i_fifo_empty           ( i_port17_in_empty ),
    .o_req0                 ( arbin17_req0 ),
    .o_req1                 ( arbin17_req1 ),
    .o_req2                 ( arbin17_req2 ),
    .i_gnt0                 ( arbin17_gnt0 ),
    .i_gnt1                 ( arbin17_gnt1 ),
    .i_gnt2                 ( arbin17_gnt2 ),
    .o_data                 ( arbin17_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i18_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port18_in_deq ), 
    .o_fifo_offset          ( o_port18_in_offset ),
    .o_fifo_eop             ( o_port18_in_eop ), 
    .i_fifo_data            ( i_port18_in_data ),
    .i_fifo_empty           ( i_port18_in_empty ),
    .o_req0                 ( arbin18_req0 ),
    .o_req1                 ( arbin18_req1 ),
    .o_req2                 ( arbin18_req2 ),
    .i_gnt0                 ( arbin18_gnt0 ),
    .i_gnt1                 ( arbin18_gnt1 ),
    .i_gnt2                 ( arbin18_gnt2 ),
    .o_data                 ( arbin18_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i19_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port19_in_deq ), 
    .o_fifo_offset          ( o_port19_in_offset ),
    .o_fifo_eop             ( o_port19_in_eop ), 
    .i_fifo_data            ( i_port19_in_data ),
    .i_fifo_empty           ( i_port19_in_empty ),
    .o_req0                 ( arbin19_req0 ),
    .o_req1                 ( arbin19_req1 ),
    .o_req2                 ( arbin19_req2 ),
    .i_gnt0                 ( arbin19_gnt0 ),
    .i_gnt1                 ( arbin19_gnt1 ),
    .i_gnt2                 ( arbin19_gnt2 ),
    .o_data                 ( arbin19_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i20_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port20_in_deq ), 
    .o_fifo_offset          ( o_port20_in_offset ),
    .o_fifo_eop             ( o_port20_in_eop ), 
    .i_fifo_data            ( i_port20_in_data ),
    .i_fifo_empty           ( i_port20_in_empty ),
    .o_req0                 ( arbin20_req0 ),
    .o_req1                 ( arbin20_req1 ),
    .o_req2                 ( arbin20_req2 ),
    .i_gnt0                 ( arbin20_gnt0 ),
    .i_gnt1                 ( arbin20_gnt1 ),
    .i_gnt2                 ( arbin20_gnt2 ),
    .o_data                 ( arbin20_data )
  );

  xbar_arb_in # (
    .ARM_MODE               ( 0 )
  ) i21_xbar_arb_in (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .i_board_id             ( i_board_id ),
    .o_fifo_deq             ( o_port21_in_deq ), 
    .o_fifo_offset          ( o_port21_in_offset ),
    .o_fifo_eop             ( o_port21_in_eop ), 
    .i_fifo_data            ( i_port21_in_data ),
    .i_fifo_empty           ( i_port21_in_empty ),
    .o_req0                 ( arbin21_req0 ),
    .o_req1                 ( arbin21_req1 ),
    .o_req2                 ( arbin21_req2 ),
    .i_gnt0                 ( arbin21_gnt0 ),
    .i_gnt1                 ( arbin21_gnt1 ),
    .i_gnt2                 ( arbin21_gnt2 ),
    .o_data                 ( arbin21_data )
  );

  
  // ==========================================================================
  // Output Arbiters
  // ==========================================================================
  xbar_arb_out i00_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port00_out_enq ),
    .o_fifo_offset          ( o_port00_out_offset ),
    .o_fifo_eop             ( o_port00_out_eop ),
    .o_fifo_data            ( o_port00_out_data ),
    .i_fifo_full            ( i_port00_out_full ),
    .i_fifo_packets_vc0     ( i_port00_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port00_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port00_out_packets_vc2 ),
    .i_req0                 ( arbout00_req0 ),
    .i_req1                 ( arbout00_req1 ),
    .i_req2                 ( arbout00_req2 ),
    .o_gnt0                 ( arbout00_gnt0 ),
    .o_gnt1                 ( arbout00_gnt1 ),
    .o_gnt2                 ( arbout00_gnt2 ),
    .o_mux_sel              ( arbout00_mux_sel ),
    .i_data                 ( arbout00_data )
  );

  xbar_arb_out i01_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port01_out_enq ),
    .o_fifo_offset          ( o_port01_out_offset ),
    .o_fifo_eop             ( o_port01_out_eop ),
    .o_fifo_data            ( o_port01_out_data ),
    .i_fifo_full            ( i_port01_out_full ),
    .i_fifo_packets_vc0     ( i_port01_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port01_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port01_out_packets_vc2 ),
    .i_req0                 ( arbout01_req0 ),
    .i_req1                 ( arbout01_req1 ),
    .i_req2                 ( arbout01_req2 ),
    .o_gnt0                 ( arbout01_gnt0 ),
    .o_gnt1                 ( arbout01_gnt1 ),
    .o_gnt2                 ( arbout01_gnt2 ),
    .o_mux_sel              ( arbout01_mux_sel ),
    .i_data                 ( arbout01_data )
  );

  xbar_arb_out i02_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port02_out_enq ),
    .o_fifo_offset          ( o_port02_out_offset ),
    .o_fifo_eop             ( o_port02_out_eop ),
    .o_fifo_data            ( o_port02_out_data ),
    .i_fifo_full            ( i_port02_out_full ),
    .i_fifo_packets_vc0     ( i_port02_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port02_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port02_out_packets_vc2 ),
    .i_req0                 ( arbout02_req0 ),
    .i_req1                 ( arbout02_req1 ),
    .i_req2                 ( arbout02_req2 ),
    .o_gnt0                 ( arbout02_gnt0 ),
    .o_gnt1                 ( arbout02_gnt1 ),
    .o_gnt2                 ( arbout02_gnt2 ),
    .o_mux_sel              ( arbout02_mux_sel ),
    .i_data                 ( arbout02_data )
  );

  xbar_arb_out i03_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port03_out_enq ),
    .o_fifo_offset          ( o_port03_out_offset ),
    .o_fifo_eop             ( o_port03_out_eop ),
    .o_fifo_data            ( o_port03_out_data ),
    .i_fifo_full            ( i_port03_out_full ),
    .i_fifo_packets_vc0     ( i_port03_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port03_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port03_out_packets_vc2 ),
    .i_req0                 ( arbout03_req0 ),
    .i_req1                 ( arbout03_req1 ),
    .i_req2                 ( arbout03_req2 ),
    .o_gnt0                 ( arbout03_gnt0 ),
    .o_gnt1                 ( arbout03_gnt1 ),
    .o_gnt2                 ( arbout03_gnt2 ),
    .o_mux_sel              ( arbout03_mux_sel ),
    .i_data                 ( arbout03_data )
  );

  xbar_arb_out i04_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port04_out_enq ),
    .o_fifo_offset          ( o_port04_out_offset ),
    .o_fifo_eop             ( o_port04_out_eop ),
    .o_fifo_data            ( o_port04_out_data ),
    .i_fifo_full            ( i_port04_out_full ),
    .i_fifo_packets_vc0     ( i_port04_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port04_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port04_out_packets_vc2 ),
    .i_req0                 ( arbout04_req0 ),
    .i_req1                 ( arbout04_req1 ),
    .i_req2                 ( arbout04_req2 ),
    .o_gnt0                 ( arbout04_gnt0 ),
    .o_gnt1                 ( arbout04_gnt1 ),
    .o_gnt2                 ( arbout04_gnt2 ),
    .o_mux_sel              ( arbout04_mux_sel ),
    .i_data                 ( arbout04_data )
  );

  xbar_arb_out i05_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port05_out_enq ),
    .o_fifo_offset          ( o_port05_out_offset ),
    .o_fifo_eop             ( o_port05_out_eop ),
    .o_fifo_data            ( o_port05_out_data ),
    .i_fifo_full            ( i_port05_out_full ),
    .i_fifo_packets_vc0     ( i_port05_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port05_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port05_out_packets_vc2 ),
    .i_req0                 ( arbout05_req0 ),
    .i_req1                 ( arbout05_req1 ),
    .i_req2                 ( arbout05_req2 ),
    .o_gnt0                 ( arbout05_gnt0 ),
    .o_gnt1                 ( arbout05_gnt1 ),
    .o_gnt2                 ( arbout05_gnt2 ),
    .o_mux_sel              ( arbout05_mux_sel ),
    .i_data                 ( arbout05_data )
  );

  xbar_arb_out i06_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port06_out_enq ),
    .o_fifo_offset          ( o_port06_out_offset ),
    .o_fifo_eop             ( o_port06_out_eop ),
    .o_fifo_data            ( o_port06_out_data ),
    .i_fifo_full            ( i_port06_out_full ),
    .i_fifo_packets_vc0     ( i_port06_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port06_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port06_out_packets_vc2 ),
    .i_req0                 ( arbout06_req0 ),
    .i_req1                 ( arbout06_req1 ),
    .i_req2                 ( arbout06_req2 ),
    .o_gnt0                 ( arbout06_gnt0 ),
    .o_gnt1                 ( arbout06_gnt1 ),
    .o_gnt2                 ( arbout06_gnt2 ),
    .o_mux_sel              ( arbout06_mux_sel ),
    .i_data                 ( arbout06_data )
  );

  xbar_arb_out i07_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port07_out_enq ),
    .o_fifo_offset          ( o_port07_out_offset ),
    .o_fifo_eop             ( o_port07_out_eop ),
    .o_fifo_data            ( o_port07_out_data ),
    .i_fifo_full            ( i_port07_out_full ),
    .i_fifo_packets_vc0     ( i_port07_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port07_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port07_out_packets_vc2 ),
    .i_req0                 ( arbout07_req0 ),
    .i_req1                 ( arbout07_req1 ),
    .i_req2                 ( arbout07_req2 ),
    .o_gnt0                 ( arbout07_gnt0 ),
    .o_gnt1                 ( arbout07_gnt1 ),
    .o_gnt2                 ( arbout07_gnt2 ),
    .o_mux_sel              ( arbout07_mux_sel ),
    .i_data                 ( arbout07_data )
  );

  xbar_arb_out i08_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port08_out_enq ),
    .o_fifo_offset          ( o_port08_out_offset ),
    .o_fifo_eop             ( o_port08_out_eop ),
    .o_fifo_data            ( o_port08_out_data ),
    .i_fifo_full            ( i_port08_out_full ),
    .i_fifo_packets_vc0     ( i_port08_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port08_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port08_out_packets_vc2 ),
    .i_req0                 ( arbout08_req0 ),
    .i_req1                 ( arbout08_req1 ),
    .i_req2                 ( arbout08_req2 ),
    .o_gnt0                 ( arbout08_gnt0 ),
    .o_gnt1                 ( arbout08_gnt1 ),
    .o_gnt2                 ( arbout08_gnt2 ),
    .o_mux_sel              ( arbout08_mux_sel ),
    .i_data                 ( arbout08_data )
  );

  xbar_arb_out i09_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port09_out_enq ),
    .o_fifo_offset          ( o_port09_out_offset ),
    .o_fifo_eop             ( o_port09_out_eop ),
    .o_fifo_data            ( o_port09_out_data ),
    .i_fifo_full            ( i_port09_out_full ),
    .i_fifo_packets_vc0     ( i_port09_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port09_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port09_out_packets_vc2 ),
    .i_req0                 ( arbout09_req0 ),
    .i_req1                 ( arbout09_req1 ),
    .i_req2                 ( arbout09_req2 ),
    .o_gnt0                 ( arbout09_gnt0 ),
    .o_gnt1                 ( arbout09_gnt1 ),
    .o_gnt2                 ( arbout09_gnt2 ),
    .o_mux_sel              ( arbout09_mux_sel ),
    .i_data                 ( arbout09_data )
  );

  xbar_arb_out i10_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port10_out_enq ),
    .o_fifo_offset          ( o_port10_out_offset ),
    .o_fifo_eop             ( o_port10_out_eop ),
    .o_fifo_data            ( o_port10_out_data ),
    .i_fifo_full            ( i_port10_out_full ),
    .i_fifo_packets_vc0     ( i_port10_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port10_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port10_out_packets_vc2 ),
    .i_req0                 ( arbout10_req0 ),
    .i_req1                 ( arbout10_req1 ),
    .i_req2                 ( arbout10_req2 ),
    .o_gnt0                 ( arbout10_gnt0 ),
    .o_gnt1                 ( arbout10_gnt1 ),
    .o_gnt2                 ( arbout10_gnt2 ),
    .o_mux_sel              ( arbout10_mux_sel ),
    .i_data                 ( arbout10_data )
  );

  xbar_arb_out i11_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port11_out_enq ),
    .o_fifo_offset          ( o_port11_out_offset ),
    .o_fifo_eop             ( o_port11_out_eop ),
    .o_fifo_data            ( o_port11_out_data ),
    .i_fifo_full            ( i_port11_out_full ),
    .i_fifo_packets_vc0     ( i_port11_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port11_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port11_out_packets_vc2 ),
    .i_req0                 ( arbout11_req0 ),
    .i_req1                 ( arbout11_req1 ),
    .i_req2                 ( arbout11_req2 ),
    .o_gnt0                 ( arbout11_gnt0 ),
    .o_gnt1                 ( arbout11_gnt1 ),
    .o_gnt2                 ( arbout11_gnt2 ),
    .o_mux_sel              ( arbout11_mux_sel ),
    .i_data                 ( arbout11_data )
  );

  xbar_arb_out i12_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port12_out_enq ),
    .o_fifo_offset          ( o_port12_out_offset ),
    .o_fifo_eop             ( o_port12_out_eop ),
    .o_fifo_data            ( o_port12_out_data ),
    .i_fifo_full            ( i_port12_out_full ),
    .i_fifo_packets_vc0     ( i_port12_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port12_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port12_out_packets_vc2 ),
    .i_req0                 ( arbout12_req0 ),
    .i_req1                 ( arbout12_req1 ),
    .i_req2                 ( arbout12_req2 ),
    .o_gnt0                 ( arbout12_gnt0 ),
    .o_gnt1                 ( arbout12_gnt1 ),
    .o_gnt2                 ( arbout12_gnt2 ),
    .o_mux_sel              ( arbout12_mux_sel ),
    .i_data                 ( arbout12_data )
  );

  xbar_arb_out i13_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port13_out_enq ),
    .o_fifo_offset          ( o_port13_out_offset ),
    .o_fifo_eop             ( o_port13_out_eop ),
    .o_fifo_data            ( o_port13_out_data ),
    .i_fifo_full            ( i_port13_out_full ),
    .i_fifo_packets_vc0     ( i_port13_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port13_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port13_out_packets_vc2 ),
    .i_req0                 ( arbout13_req0 ),
    .i_req1                 ( arbout13_req1 ),
    .i_req2                 ( arbout13_req2 ),
    .o_gnt0                 ( arbout13_gnt0 ),
    .o_gnt1                 ( arbout13_gnt1 ),
    .o_gnt2                 ( arbout13_gnt2 ),
    .o_mux_sel              ( arbout13_mux_sel ),
    .i_data                 ( arbout13_data )
  );

  xbar_arb_out i14_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port14_out_enq ),
    .o_fifo_offset          ( o_port14_out_offset ),
    .o_fifo_eop             ( o_port14_out_eop ),
    .o_fifo_data            ( o_port14_out_data ),
    .i_fifo_full            ( i_port14_out_full ),
    .i_fifo_packets_vc0     ( i_port14_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port14_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port14_out_packets_vc2 ),
    .i_req0                 ( arbout14_req0 ),
    .i_req1                 ( arbout14_req1 ),
    .i_req2                 ( arbout14_req2 ),
    .o_gnt0                 ( arbout14_gnt0 ),
    .o_gnt1                 ( arbout14_gnt1 ),
    .o_gnt2                 ( arbout14_gnt2 ),
    .o_mux_sel              ( arbout14_mux_sel ),
    .i_data                 ( arbout14_data )
  );

  xbar_arb_out i15_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port15_out_enq ),
    .o_fifo_offset          ( o_port15_out_offset ),
    .o_fifo_eop             ( o_port15_out_eop ),
    .o_fifo_data            ( o_port15_out_data ),
    .i_fifo_full            ( i_port15_out_full ),
    .i_fifo_packets_vc0     ( i_port15_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port15_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port15_out_packets_vc2 ),
    .i_req0                 ( arbout15_req0 ),
    .i_req1                 ( arbout15_req1 ),
    .i_req2                 ( arbout15_req2 ),
    .o_gnt0                 ( arbout15_gnt0 ),
    .o_gnt1                 ( arbout15_gnt1 ),
    .o_gnt2                 ( arbout15_gnt2 ),
    .o_mux_sel              ( arbout15_mux_sel ),
    .i_data                 ( arbout15_data )
  );

  xbar_arb_out i16_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port16_out_enq ),
    .o_fifo_offset          ( o_port16_out_offset ),
    .o_fifo_eop             ( o_port16_out_eop ),
    .o_fifo_data            ( o_port16_out_data ),
    .i_fifo_full            ( i_port16_out_full ),
    .i_fifo_packets_vc0     ( i_port16_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port16_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port16_out_packets_vc2 ),
    .i_req0                 ( arbout16_req0 ),
    .i_req1                 ( arbout16_req1 ),
    .i_req2                 ( arbout16_req2 ),
    .o_gnt0                 ( arbout16_gnt0 ),
    .o_gnt1                 ( arbout16_gnt1 ),
    .o_gnt2                 ( arbout16_gnt2 ),
    .o_mux_sel              ( arbout16_mux_sel ),
    .i_data                 ( arbout16_data )
  );

  xbar_arb_out i17_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port17_out_enq ),
    .o_fifo_offset          ( o_port17_out_offset ),
    .o_fifo_eop             ( o_port17_out_eop ),
    .o_fifo_data            ( o_port17_out_data ),
    .i_fifo_full            ( i_port17_out_full ),
    .i_fifo_packets_vc0     ( i_port17_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port17_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port17_out_packets_vc2 ),
    .i_req0                 ( arbout17_req0 ),
    .i_req1                 ( arbout17_req1 ),
    .i_req2                 ( arbout17_req2 ),
    .o_gnt0                 ( arbout17_gnt0 ),
    .o_gnt1                 ( arbout17_gnt1 ),
    .o_gnt2                 ( arbout17_gnt2 ),
    .o_mux_sel              ( arbout17_mux_sel ),
    .i_data                 ( arbout17_data )
  );

  xbar_arb_out i18_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port18_out_enq ),
    .o_fifo_offset          ( o_port18_out_offset ),
    .o_fifo_eop             ( o_port18_out_eop ),
    .o_fifo_data            ( o_port18_out_data ),
    .i_fifo_full            ( i_port18_out_full ),
    .i_fifo_packets_vc0     ( i_port18_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port18_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port18_out_packets_vc2 ),
    .i_req0                 ( arbout18_req0 ),
    .i_req1                 ( arbout18_req1 ),
    .i_req2                 ( arbout18_req2 ),
    .o_gnt0                 ( arbout18_gnt0 ),
    .o_gnt1                 ( arbout18_gnt1 ),
    .o_gnt2                 ( arbout18_gnt2 ),
    .o_mux_sel              ( arbout18_mux_sel ),
    .i_data                 ( arbout18_data )
  );

  xbar_arb_out i19_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port19_out_enq ),
    .o_fifo_offset          ( o_port19_out_offset ),
    .o_fifo_eop             ( o_port19_out_eop ),
    .o_fifo_data            ( o_port19_out_data ),
    .i_fifo_full            ( i_port19_out_full ),
    .i_fifo_packets_vc0     ( i_port19_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port19_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port19_out_packets_vc2 ),
    .i_req0                 ( arbout19_req0 ),
    .i_req1                 ( arbout19_req1 ),
    .i_req2                 ( arbout19_req2 ),
    .o_gnt0                 ( arbout19_gnt0 ),
    .o_gnt1                 ( arbout19_gnt1 ),
    .o_gnt2                 ( arbout19_gnt2 ),
    .o_mux_sel              ( arbout19_mux_sel ),
    .i_data                 ( arbout19_data )
  );

  xbar_arb_out i20_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port20_out_enq ),
    .o_fifo_offset          ( o_port20_out_offset ),
    .o_fifo_eop             ( o_port20_out_eop ),
    .o_fifo_data            ( o_port20_out_data ),
    .i_fifo_full            ( i_port20_out_full ),
    .i_fifo_packets_vc0     ( i_port20_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port20_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port20_out_packets_vc2 ),
    .i_req0                 ( arbout20_req0 ),
    .i_req1                 ( arbout20_req1 ),
    .i_req2                 ( arbout20_req2 ),
    .o_gnt0                 ( arbout20_gnt0 ),
    .o_gnt1                 ( arbout20_gnt1 ),
    .o_gnt2                 ( arbout20_gnt2 ),
    .o_mux_sel              ( arbout20_mux_sel ),
    .i_data                 ( arbout20_data )
  );

  xbar_arb_out i21_xbar_arb_out (
    .clk                    ( clk_xbar ),
    .rst                    ( rst_xbar ),
    .o_fifo_enq             ( o_port21_out_enq ),
    .o_fifo_offset          ( o_port21_out_offset ),
    .o_fifo_eop             ( o_port21_out_eop ),
    .o_fifo_data            ( o_port21_out_data ),
    .i_fifo_full            ( i_port21_out_full ),
    .i_fifo_packets_vc0     ( i_port21_out_packets_vc0 ),
    .i_fifo_packets_vc1     ( i_port21_out_packets_vc1 ),
    .i_fifo_packets_vc2     ( i_port21_out_packets_vc2 ),
    .i_req0                 ( arbout21_req0 ),
    .i_req1                 ( arbout21_req1 ),
    .i_req2                 ( arbout21_req2 ),
    .o_gnt0                 ( arbout21_gnt0 ),
    .o_gnt1                 ( arbout21_gnt1 ),
    .o_gnt2                 ( arbout21_gnt2 ),
    .o_mux_sel              ( arbout21_mux_sel ),
    .i_data                 ( arbout21_data )
  );



  // ==========================================================================
  // Switching fabric: Data muxes
  // ==========================================================================
  xbar_mux i00_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout00_mux_sel ),
    .o_data                 ( arbout00_data )
  );

  xbar_mux i01_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout01_mux_sel ),
    .o_data                 ( arbout01_data )
  );

  xbar_mux i02_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout02_mux_sel ),
    .o_data                 ( arbout02_data )
  );

  xbar_mux i03_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout03_mux_sel ),
    .o_data                 ( arbout03_data )
  );

  xbar_mux i04_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout04_mux_sel ),
    .o_data                 ( arbout04_data )
  );

  xbar_mux i05_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout05_mux_sel ),
    .o_data                 ( arbout05_data )
  );

  xbar_mux i06_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout06_mux_sel ),
    .o_data                 ( arbout06_data )
  );

  xbar_mux i07_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout07_mux_sel ),
    .o_data                 ( arbout07_data )
  );

  xbar_mux i08_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout08_mux_sel ),
    .o_data                 ( arbout08_data )
  );

  xbar_mux i09_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout09_mux_sel ),
    .o_data                 ( arbout09_data )
  );

  xbar_mux i10_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout10_mux_sel ),
    .o_data                 ( arbout10_data )
  );

  xbar_mux i11_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout11_mux_sel ),
    .o_data                 ( arbout11_data )
  );

  xbar_mux i12_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout12_mux_sel ),
    .o_data                 ( arbout12_data )
  );

  xbar_mux i13_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout13_mux_sel ),
    .o_data                 ( arbout13_data )
  );

  xbar_mux i14_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout14_mux_sel ),
    .o_data                 ( arbout14_data )
  );

  xbar_mux i15_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout15_mux_sel ),
    .o_data                 ( arbout15_data )
  );

  xbar_mux i16_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout16_mux_sel ),
    .o_data                 ( arbout16_data )
  );

  xbar_mux i17_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout17_mux_sel ),
    .o_data                 ( arbout17_data )
  );

  xbar_mux i18_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout18_mux_sel ),
    .o_data                 ( arbout18_data )
  );

  xbar_mux i19_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout19_mux_sel ),
    .o_data                 ( arbout19_data )
  );

  xbar_mux i20_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout20_mux_sel ),
    .o_data                 ( arbout20_data )
  );

  xbar_mux i21_xbar_mux (
    .clk                    ( clk_xbar ),
    .i_data00               ( arbin00_data ),
    .i_data01               ( arbin01_data ),
    .i_data02               ( arbin02_data ),
    .i_data03               ( arbin03_data ),
    .i_data04               ( arbin04_data ),
    .i_data05               ( arbin05_data ),
    .i_data06               ( arbin06_data ),
    .i_data07               ( arbin07_data ),
    .i_data08               ( arbin08_data ),
    .i_data09               ( arbin09_data ),
    .i_data10               ( arbin10_data ),
    .i_data11               ( arbin11_data ),
    .i_data12               ( arbin12_data ),
    .i_data13               ( arbin13_data ),
    .i_data14               ( arbin14_data ),
    .i_data15               ( arbin15_data ),
    .i_data16               ( arbin16_data ),
    .i_data17               ( arbin17_data ),
    .i_data18               ( arbin18_data ),
    .i_data19               ( arbin19_data ),
    .i_data20               ( arbin20_data ),
    .i_data21               ( arbin21_data ),
    .i_sel                  ( arbout21_mux_sel ),
    .o_data                 ( arbout21_data )
  );

  
  // ==========================================================================
  // Request stiching
  // ==========================================================================
  assign arbout00_req0 = {
    arbin21_req0[0], arbin20_req0[0], arbin19_req0[0], arbin18_req0[0],
    arbin17_req0[0], arbin16_req0[0], arbin15_req0[0], arbin14_req0[0],
    arbin13_req0[0], arbin12_req0[0], arbin11_req0[0], arbin10_req0[0],
    arbin09_req0[0], arbin08_req0[0], arbin07_req0[0], arbin06_req0[0],
    arbin05_req0[0], arbin04_req0[0], arbin03_req0[0], arbin02_req0[0],
    arbin01_req0[0], arbin00_req0[0]};

  assign arbout01_req0 = {
    arbin21_req0[1], arbin20_req0[1], arbin19_req0[1], arbin18_req0[1],
    arbin17_req0[1], arbin16_req0[1], arbin15_req0[1], arbin14_req0[1],
    arbin13_req0[1], arbin12_req0[1], arbin11_req0[1], arbin10_req0[1],
    arbin09_req0[1], arbin08_req0[1], arbin07_req0[1], arbin06_req0[1],
    arbin05_req0[1], arbin04_req0[1], arbin03_req0[1], arbin02_req0[1],
    arbin01_req0[1], arbin00_req0[1]};

  assign arbout02_req0 = {
    arbin21_req0[2], arbin20_req0[2], arbin19_req0[2], arbin18_req0[2],
    arbin17_req0[2], arbin16_req0[2], arbin15_req0[2], arbin14_req0[2],
    arbin13_req0[2], arbin12_req0[2], arbin11_req0[2], arbin10_req0[2],
    arbin09_req0[2], arbin08_req0[2], arbin07_req0[2], arbin06_req0[2],
    arbin05_req0[2], arbin04_req0[2], arbin03_req0[2], arbin02_req0[2],
    arbin01_req0[2], arbin00_req0[2]};

  assign arbout03_req0 = {
    arbin21_req0[3], arbin20_req0[3], arbin19_req0[3], arbin18_req0[3],
    arbin17_req0[3], arbin16_req0[3], arbin15_req0[3], arbin14_req0[3],
    arbin13_req0[3], arbin12_req0[3], arbin11_req0[3], arbin10_req0[3],
    arbin09_req0[3], arbin08_req0[3], arbin07_req0[3], arbin06_req0[3],
    arbin05_req0[3], arbin04_req0[3], arbin03_req0[3], arbin02_req0[3],
    arbin01_req0[3], arbin00_req0[3]};

  assign arbout04_req0 = {
    arbin21_req0[4], arbin20_req0[4], arbin19_req0[4], arbin18_req0[4],
    arbin17_req0[4], arbin16_req0[4], arbin15_req0[4], arbin14_req0[4],
    arbin13_req0[4], arbin12_req0[4], arbin11_req0[4], arbin10_req0[4],
    arbin09_req0[4], arbin08_req0[4], arbin07_req0[4], arbin06_req0[4],
    arbin05_req0[4], arbin04_req0[4], arbin03_req0[4], arbin02_req0[4],
    arbin01_req0[4], arbin00_req0[4]};

  assign arbout05_req0 = {
    arbin21_req0[5], arbin20_req0[5], arbin19_req0[5], arbin18_req0[5],
    arbin17_req0[5], arbin16_req0[5], arbin15_req0[5], arbin14_req0[5],
    arbin13_req0[5], arbin12_req0[5], arbin11_req0[5], arbin10_req0[5],
    arbin09_req0[5], arbin08_req0[5], arbin07_req0[5], arbin06_req0[5],
    arbin05_req0[5], arbin04_req0[5], arbin03_req0[5], arbin02_req0[5],
    arbin01_req0[5], arbin00_req0[5]};

  assign arbout06_req0 = {
    arbin21_req0[6], arbin20_req0[6], arbin19_req0[6], arbin18_req0[6],
    arbin17_req0[6], arbin16_req0[6], arbin15_req0[6], arbin14_req0[6],
    arbin13_req0[6], arbin12_req0[6], arbin11_req0[6], arbin10_req0[6],
    arbin09_req0[6], arbin08_req0[6], arbin07_req0[6], arbin06_req0[6],
    arbin05_req0[6], arbin04_req0[6], arbin03_req0[6], arbin02_req0[6],
    arbin01_req0[6], arbin00_req0[6]};

  assign arbout07_req0 = {
    arbin21_req0[7], arbin20_req0[7], arbin19_req0[7], arbin18_req0[7],
    arbin17_req0[7], arbin16_req0[7], arbin15_req0[7], arbin14_req0[7],
    arbin13_req0[7], arbin12_req0[7], arbin11_req0[7], arbin10_req0[7],
    arbin09_req0[7], arbin08_req0[7], arbin07_req0[7], arbin06_req0[7],
    arbin05_req0[7], arbin04_req0[7], arbin03_req0[7], arbin02_req0[7],
    arbin01_req0[7], arbin00_req0[7]};

  assign arbout08_req0 = {
    arbin21_req0[8], arbin20_req0[8], arbin19_req0[8], arbin18_req0[8],
    arbin17_req0[8], arbin16_req0[8], arbin15_req0[8], arbin14_req0[8],
    arbin13_req0[8], arbin12_req0[8], arbin11_req0[8], arbin10_req0[8],
    arbin09_req0[8], arbin08_req0[8], arbin07_req0[8], arbin06_req0[8],
    arbin05_req0[8], arbin04_req0[8], arbin03_req0[8], arbin02_req0[8],
    arbin01_req0[8], arbin00_req0[8]};

  assign arbout09_req0 = {
    arbin21_req0[9], arbin20_req0[9], arbin19_req0[9], arbin18_req0[9],
    arbin17_req0[9], arbin16_req0[9], arbin15_req0[9], arbin14_req0[9],
    arbin13_req0[9], arbin12_req0[9], arbin11_req0[9], arbin10_req0[9],
    arbin09_req0[9], arbin08_req0[9], arbin07_req0[9], arbin06_req0[9],
    arbin05_req0[9], arbin04_req0[9], arbin03_req0[9], arbin02_req0[9],
    arbin01_req0[9], arbin00_req0[9]};

  assign arbout10_req0 = {
    arbin21_req0[10], arbin20_req0[10], arbin19_req0[10], arbin18_req0[10],
    arbin17_req0[10], arbin16_req0[10], arbin15_req0[10], arbin14_req0[10],
    arbin13_req0[10], arbin12_req0[10], arbin11_req0[10], arbin10_req0[10],
    arbin09_req0[10], arbin08_req0[10], arbin07_req0[10], arbin06_req0[10],
    arbin05_req0[10], arbin04_req0[10], arbin03_req0[10], arbin02_req0[10],
    arbin01_req0[10], arbin00_req0[10]};

  assign arbout11_req0 = {
    arbin21_req0[11], arbin20_req0[11], arbin19_req0[11], arbin18_req0[11],
    arbin17_req0[11], arbin16_req0[11], arbin15_req0[11], arbin14_req0[11],
    arbin13_req0[11], arbin12_req0[11], arbin11_req0[11], arbin10_req0[11],
    arbin09_req0[11], arbin08_req0[11], arbin07_req0[11], arbin06_req0[11],
    arbin05_req0[11], arbin04_req0[11], arbin03_req0[11], arbin02_req0[11],
    arbin01_req0[11], arbin00_req0[11]};

  assign arbout12_req0 = {
    arbin21_req0[12], arbin20_req0[12], arbin19_req0[12], arbin18_req0[12],
    arbin17_req0[12], arbin16_req0[12], arbin15_req0[12], arbin14_req0[12],
    arbin13_req0[12], arbin12_req0[12], arbin11_req0[12], arbin10_req0[12],
    arbin09_req0[12], arbin08_req0[12], arbin07_req0[12], arbin06_req0[12],
    arbin05_req0[12], arbin04_req0[12], arbin03_req0[12], arbin02_req0[12],
    arbin01_req0[12], arbin00_req0[12]};

  assign arbout13_req0 = {
    arbin21_req0[13], arbin20_req0[13], arbin19_req0[13], arbin18_req0[13],
    arbin17_req0[13], arbin16_req0[13], arbin15_req0[13], arbin14_req0[13],
    arbin13_req0[13], arbin12_req0[13], arbin11_req0[13], arbin10_req0[13],
    arbin09_req0[13], arbin08_req0[13], arbin07_req0[13], arbin06_req0[13],
    arbin05_req0[13], arbin04_req0[13], arbin03_req0[13], arbin02_req0[13],
    arbin01_req0[13], arbin00_req0[13]};

  assign arbout14_req0 = {
    arbin21_req0[14], arbin20_req0[14], arbin19_req0[14], arbin18_req0[14],
    arbin17_req0[14], arbin16_req0[14], arbin15_req0[14], arbin14_req0[14],
    arbin13_req0[14], arbin12_req0[14], arbin11_req0[14], arbin10_req0[14],
    arbin09_req0[14], arbin08_req0[14], arbin07_req0[14], arbin06_req0[14],
    arbin05_req0[14], arbin04_req0[14], arbin03_req0[14], arbin02_req0[14],
    arbin01_req0[14], arbin00_req0[14]};

  assign arbout15_req0 = {
    arbin21_req0[15], arbin20_req0[15], arbin19_req0[15], arbin18_req0[15],
    arbin17_req0[15], arbin16_req0[15], arbin15_req0[15], arbin14_req0[15],
    arbin13_req0[15], arbin12_req0[15], arbin11_req0[15], arbin10_req0[15],
    arbin09_req0[15], arbin08_req0[15], arbin07_req0[15], arbin06_req0[15],
    arbin05_req0[15], arbin04_req0[15], arbin03_req0[15], arbin02_req0[15],
    arbin01_req0[15], arbin00_req0[15]};

  assign arbout16_req0 = {
    arbin21_req0[16], arbin20_req0[16], arbin19_req0[16], arbin18_req0[16],
    arbin17_req0[16], arbin16_req0[16], arbin15_req0[16], arbin14_req0[16],
    arbin13_req0[16], arbin12_req0[16], arbin11_req0[16], arbin10_req0[16],
    arbin09_req0[16], arbin08_req0[16], arbin07_req0[16], arbin06_req0[16],
    arbin05_req0[16], arbin04_req0[16], arbin03_req0[16], arbin02_req0[16],
    arbin01_req0[16], arbin00_req0[16]};

  assign arbout17_req0 = {
    arbin21_req0[17], arbin20_req0[17], arbin19_req0[17], arbin18_req0[17],
    arbin17_req0[17], arbin16_req0[17], arbin15_req0[17], arbin14_req0[17],
    arbin13_req0[17], arbin12_req0[17], arbin11_req0[17], arbin10_req0[17],
    arbin09_req0[17], arbin08_req0[17], arbin07_req0[17], arbin06_req0[17],
    arbin05_req0[17], arbin04_req0[17], arbin03_req0[17], arbin02_req0[17],
    arbin01_req0[17], arbin00_req0[17]};

  assign arbout18_req0 = {
    arbin21_req0[18], arbin20_req0[18], arbin19_req0[18], arbin18_req0[18],
    arbin17_req0[18], arbin16_req0[18], arbin15_req0[18], arbin14_req0[18],
    arbin13_req0[18], arbin12_req0[18], arbin11_req0[18], arbin10_req0[18],
    arbin09_req0[18], arbin08_req0[18], arbin07_req0[18], arbin06_req0[18],
    arbin05_req0[18], arbin04_req0[18], arbin03_req0[18], arbin02_req0[18],
    arbin01_req0[18], arbin00_req0[18]};

  assign arbout19_req0 = {
    arbin21_req0[19], arbin20_req0[19], arbin19_req0[19], arbin18_req0[19],
    arbin17_req0[19], arbin16_req0[19], arbin15_req0[19], arbin14_req0[19],
    arbin13_req0[19], arbin12_req0[19], arbin11_req0[19], arbin10_req0[19],
    arbin09_req0[19], arbin08_req0[19], arbin07_req0[19], arbin06_req0[19],
    arbin05_req0[19], arbin04_req0[19], arbin03_req0[19], arbin02_req0[19],
    arbin01_req0[19], arbin00_req0[19]};

  assign arbout20_req0 = {
    arbin21_req0[20], arbin20_req0[20], arbin19_req0[20], arbin18_req0[20],
    arbin17_req0[20], arbin16_req0[20], arbin15_req0[20], arbin14_req0[20],
    arbin13_req0[20], arbin12_req0[20], arbin11_req0[20], arbin10_req0[20],
    arbin09_req0[20], arbin08_req0[20], arbin07_req0[20], arbin06_req0[20],
    arbin05_req0[20], arbin04_req0[20], arbin03_req0[20], arbin02_req0[20],
    arbin01_req0[20], arbin00_req0[20]};

  assign arbout21_req0 = {
    arbin21_req0[21], arbin20_req0[21], arbin19_req0[21], arbin18_req0[21],
    arbin17_req0[21], arbin16_req0[21], arbin15_req0[21], arbin14_req0[21],
    arbin13_req0[21], arbin12_req0[21], arbin11_req0[21], arbin10_req0[21],
    arbin09_req0[21], arbin08_req0[21], arbin07_req0[21], arbin06_req0[21],
    arbin05_req0[21], arbin04_req0[21], arbin03_req0[21], arbin02_req0[21],
    arbin01_req0[21], arbin00_req0[21]};

  assign arbout00_req1 = {
    arbin21_req1[0], arbin20_req1[0], arbin19_req1[0], arbin18_req1[0],
    arbin17_req1[0], arbin16_req1[0], arbin15_req1[0], arbin14_req1[0],
    arbin13_req1[0], arbin12_req1[0], arbin11_req1[0], arbin10_req1[0],
    arbin09_req1[0], arbin08_req1[0], arbin07_req1[0], arbin06_req1[0],
    arbin05_req1[0], arbin04_req1[0], arbin03_req1[0], arbin02_req1[0],
    arbin01_req1[0], arbin00_req1[0]};

  assign arbout01_req1 = {
    arbin21_req1[1], arbin20_req1[1], arbin19_req1[1], arbin18_req1[1],
    arbin17_req1[1], arbin16_req1[1], arbin15_req1[1], arbin14_req1[1],
    arbin13_req1[1], arbin12_req1[1], arbin11_req1[1], arbin10_req1[1],
    arbin09_req1[1], arbin08_req1[1], arbin07_req1[1], arbin06_req1[1],
    arbin05_req1[1], arbin04_req1[1], arbin03_req1[1], arbin02_req1[1],
    arbin01_req1[1], arbin00_req1[1]};

  assign arbout02_req1 = {
    arbin21_req1[2], arbin20_req1[2], arbin19_req1[2], arbin18_req1[2],
    arbin17_req1[2], arbin16_req1[2], arbin15_req1[2], arbin14_req1[2],
    arbin13_req1[2], arbin12_req1[2], arbin11_req1[2], arbin10_req1[2],
    arbin09_req1[2], arbin08_req1[2], arbin07_req1[2], arbin06_req1[2],
    arbin05_req1[2], arbin04_req1[2], arbin03_req1[2], arbin02_req1[2],
    arbin01_req1[2], arbin00_req1[2]};

  assign arbout03_req1 = {
    arbin21_req1[3], arbin20_req1[3], arbin19_req1[3], arbin18_req1[3],
    arbin17_req1[3], arbin16_req1[3], arbin15_req1[3], arbin14_req1[3],
    arbin13_req1[3], arbin12_req1[3], arbin11_req1[3], arbin10_req1[3],
    arbin09_req1[3], arbin08_req1[3], arbin07_req1[3], arbin06_req1[3],
    arbin05_req1[3], arbin04_req1[3], arbin03_req1[3], arbin02_req1[3],
    arbin01_req1[3], arbin00_req1[3]};

  assign arbout04_req1 = {
    arbin21_req1[4], arbin20_req1[4], arbin19_req1[4], arbin18_req1[4],
    arbin17_req1[4], arbin16_req1[4], arbin15_req1[4], arbin14_req1[4],
    arbin13_req1[4], arbin12_req1[4], arbin11_req1[4], arbin10_req1[4],
    arbin09_req1[4], arbin08_req1[4], arbin07_req1[4], arbin06_req1[4],
    arbin05_req1[4], arbin04_req1[4], arbin03_req1[4], arbin02_req1[4],
    arbin01_req1[4], arbin00_req1[4]};

  assign arbout05_req1 = {
    arbin21_req1[5], arbin20_req1[5], arbin19_req1[5], arbin18_req1[5],
    arbin17_req1[5], arbin16_req1[5], arbin15_req1[5], arbin14_req1[5],
    arbin13_req1[5], arbin12_req1[5], arbin11_req1[5], arbin10_req1[5],
    arbin09_req1[5], arbin08_req1[5], arbin07_req1[5], arbin06_req1[5],
    arbin05_req1[5], arbin04_req1[5], arbin03_req1[5], arbin02_req1[5],
    arbin01_req1[5], arbin00_req1[5]};

  assign arbout06_req1 = {
    arbin21_req1[6], arbin20_req1[6], arbin19_req1[6], arbin18_req1[6],
    arbin17_req1[6], arbin16_req1[6], arbin15_req1[6], arbin14_req1[6],
    arbin13_req1[6], arbin12_req1[6], arbin11_req1[6], arbin10_req1[6],
    arbin09_req1[6], arbin08_req1[6], arbin07_req1[6], arbin06_req1[6],
    arbin05_req1[6], arbin04_req1[6], arbin03_req1[6], arbin02_req1[6],
    arbin01_req1[6], arbin00_req1[6]};

  assign arbout07_req1 = {
    arbin21_req1[7], arbin20_req1[7], arbin19_req1[7], arbin18_req1[7],
    arbin17_req1[7], arbin16_req1[7], arbin15_req1[7], arbin14_req1[7],
    arbin13_req1[7], arbin12_req1[7], arbin11_req1[7], arbin10_req1[7],
    arbin09_req1[7], arbin08_req1[7], arbin07_req1[7], arbin06_req1[7],
    arbin05_req1[7], arbin04_req1[7], arbin03_req1[7], arbin02_req1[7],
    arbin01_req1[7], arbin00_req1[7]};

  assign arbout08_req1 = {
    arbin21_req1[8], arbin20_req1[8], arbin19_req1[8], arbin18_req1[8],
    arbin17_req1[8], arbin16_req1[8], arbin15_req1[8], arbin14_req1[8],
    arbin13_req1[8], arbin12_req1[8], arbin11_req1[8], arbin10_req1[8],
    arbin09_req1[8], arbin08_req1[8], arbin07_req1[8], arbin06_req1[8],
    arbin05_req1[8], arbin04_req1[8], arbin03_req1[8], arbin02_req1[8],
    arbin01_req1[8], arbin00_req1[8]};

  assign arbout09_req1 = {
    arbin21_req1[9], arbin20_req1[9], arbin19_req1[9], arbin18_req1[9],
    arbin17_req1[9], arbin16_req1[9], arbin15_req1[9], arbin14_req1[9],
    arbin13_req1[9], arbin12_req1[9], arbin11_req1[9], arbin10_req1[9],
    arbin09_req1[9], arbin08_req1[9], arbin07_req1[9], arbin06_req1[9],
    arbin05_req1[9], arbin04_req1[9], arbin03_req1[9], arbin02_req1[9],
    arbin01_req1[9], arbin00_req1[9]};

  assign arbout10_req1 = {
    arbin21_req1[10], arbin20_req1[10], arbin19_req1[10], arbin18_req1[10],
    arbin17_req1[10], arbin16_req1[10], arbin15_req1[10], arbin14_req1[10],
    arbin13_req1[10], arbin12_req1[10], arbin11_req1[10], arbin10_req1[10],
    arbin09_req1[10], arbin08_req1[10], arbin07_req1[10], arbin06_req1[10],
    arbin05_req1[10], arbin04_req1[10], arbin03_req1[10], arbin02_req1[10],
    arbin01_req1[10], arbin00_req1[10]};

  assign arbout11_req1 = {
    arbin21_req1[11], arbin20_req1[11], arbin19_req1[11], arbin18_req1[11],
    arbin17_req1[11], arbin16_req1[11], arbin15_req1[11], arbin14_req1[11],
    arbin13_req1[11], arbin12_req1[11], arbin11_req1[11], arbin10_req1[11],
    arbin09_req1[11], arbin08_req1[11], arbin07_req1[11], arbin06_req1[11],
    arbin05_req1[11], arbin04_req1[11], arbin03_req1[11], arbin02_req1[11],
    arbin01_req1[11], arbin00_req1[11]};

  assign arbout12_req1 = {
    arbin21_req1[12], arbin20_req1[12], arbin19_req1[12], arbin18_req1[12],
    arbin17_req1[12], arbin16_req1[12], arbin15_req1[12], arbin14_req1[12],
    arbin13_req1[12], arbin12_req1[12], arbin11_req1[12], arbin10_req1[12],
    arbin09_req1[12], arbin08_req1[12], arbin07_req1[12], arbin06_req1[12],
    arbin05_req1[12], arbin04_req1[12], arbin03_req1[12], arbin02_req1[12],
    arbin01_req1[12], arbin00_req1[12]};

  assign arbout13_req1 = {
    arbin21_req1[13], arbin20_req1[13], arbin19_req1[13], arbin18_req1[13],
    arbin17_req1[13], arbin16_req1[13], arbin15_req1[13], arbin14_req1[13],
    arbin13_req1[13], arbin12_req1[13], arbin11_req1[13], arbin10_req1[13],
    arbin09_req1[13], arbin08_req1[13], arbin07_req1[13], arbin06_req1[13],
    arbin05_req1[13], arbin04_req1[13], arbin03_req1[13], arbin02_req1[13],
    arbin01_req1[13], arbin00_req1[13]};

  assign arbout14_req1 = {
    arbin21_req1[14], arbin20_req1[14], arbin19_req1[14], arbin18_req1[14],
    arbin17_req1[14], arbin16_req1[14], arbin15_req1[14], arbin14_req1[14],
    arbin13_req1[14], arbin12_req1[14], arbin11_req1[14], arbin10_req1[14],
    arbin09_req1[14], arbin08_req1[14], arbin07_req1[14], arbin06_req1[14],
    arbin05_req1[14], arbin04_req1[14], arbin03_req1[14], arbin02_req1[14],
    arbin01_req1[14], arbin00_req1[14]};

  assign arbout15_req1 = {
    arbin21_req1[15], arbin20_req1[15], arbin19_req1[15], arbin18_req1[15],
    arbin17_req1[15], arbin16_req1[15], arbin15_req1[15], arbin14_req1[15],
    arbin13_req1[15], arbin12_req1[15], arbin11_req1[15], arbin10_req1[15],
    arbin09_req1[15], arbin08_req1[15], arbin07_req1[15], arbin06_req1[15],
    arbin05_req1[15], arbin04_req1[15], arbin03_req1[15], arbin02_req1[15],
    arbin01_req1[15], arbin00_req1[15]};

  assign arbout16_req1 = {
    arbin21_req1[16], arbin20_req1[16], arbin19_req1[16], arbin18_req1[16],
    arbin17_req1[16], arbin16_req1[16], arbin15_req1[16], arbin14_req1[16],
    arbin13_req1[16], arbin12_req1[16], arbin11_req1[16], arbin10_req1[16],
    arbin09_req1[16], arbin08_req1[16], arbin07_req1[16], arbin06_req1[16],
    arbin05_req1[16], arbin04_req1[16], arbin03_req1[16], arbin02_req1[16],
    arbin01_req1[16], arbin00_req1[16]};

  assign arbout17_req1 = {
    arbin21_req1[17], arbin20_req1[17], arbin19_req1[17], arbin18_req1[17],
    arbin17_req1[17], arbin16_req1[17], arbin15_req1[17], arbin14_req1[17],
    arbin13_req1[17], arbin12_req1[17], arbin11_req1[17], arbin10_req1[17],
    arbin09_req1[17], arbin08_req1[17], arbin07_req1[17], arbin06_req1[17],
    arbin05_req1[17], arbin04_req1[17], arbin03_req1[17], arbin02_req1[17],
    arbin01_req1[17], arbin00_req1[17]};

  assign arbout18_req1 = {
    arbin21_req1[18], arbin20_req1[18], arbin19_req1[18], arbin18_req1[18],
    arbin17_req1[18], arbin16_req1[18], arbin15_req1[18], arbin14_req1[18],
    arbin13_req1[18], arbin12_req1[18], arbin11_req1[18], arbin10_req1[18],
    arbin09_req1[18], arbin08_req1[18], arbin07_req1[18], arbin06_req1[18],
    arbin05_req1[18], arbin04_req1[18], arbin03_req1[18], arbin02_req1[18],
    arbin01_req1[18], arbin00_req1[18]};

  assign arbout19_req1 = {
    arbin21_req1[19], arbin20_req1[19], arbin19_req1[19], arbin18_req1[19],
    arbin17_req1[19], arbin16_req1[19], arbin15_req1[19], arbin14_req1[19],
    arbin13_req1[19], arbin12_req1[19], arbin11_req1[19], arbin10_req1[19],
    arbin09_req1[19], arbin08_req1[19], arbin07_req1[19], arbin06_req1[19],
    arbin05_req1[19], arbin04_req1[19], arbin03_req1[19], arbin02_req1[19],
    arbin01_req1[19], arbin00_req1[19]};

  assign arbout20_req1 = {
    arbin21_req1[20], arbin20_req1[20], arbin19_req1[20], arbin18_req1[20],
    arbin17_req1[20], arbin16_req1[20], arbin15_req1[20], arbin14_req1[20],
    arbin13_req1[20], arbin12_req1[20], arbin11_req1[20], arbin10_req1[20],
    arbin09_req1[20], arbin08_req1[20], arbin07_req1[20], arbin06_req1[20],
    arbin05_req1[20], arbin04_req1[20], arbin03_req1[20], arbin02_req1[20],
    arbin01_req1[20], arbin00_req1[20]};

  assign arbout21_req1 = {
    arbin21_req1[21], arbin20_req1[21], arbin19_req1[21], arbin18_req1[21],
    arbin17_req1[21], arbin16_req1[21], arbin15_req1[21], arbin14_req1[21],
    arbin13_req1[21], arbin12_req1[21], arbin11_req1[21], arbin10_req1[21],
    arbin09_req1[21], arbin08_req1[21], arbin07_req1[21], arbin06_req1[21],
    arbin05_req1[21], arbin04_req1[21], arbin03_req1[21], arbin02_req1[21],
    arbin01_req1[21], arbin00_req1[21]};

  assign arbout00_req2 = {
    arbin21_req2[0], arbin20_req2[0], arbin19_req2[0], arbin18_req2[0],
    arbin17_req2[0], arbin16_req2[0], arbin15_req2[0], arbin14_req2[0],
    arbin13_req2[0], arbin12_req2[0], arbin11_req2[0], arbin10_req2[0],
    arbin09_req2[0], arbin08_req2[0], arbin07_req2[0], arbin06_req2[0],
    arbin05_req2[0], arbin04_req2[0], arbin03_req2[0], arbin02_req2[0],
    arbin01_req2[0], arbin00_req2[0]};

  assign arbout01_req2 = {
    arbin21_req2[1], arbin20_req2[1], arbin19_req2[1], arbin18_req2[1],
    arbin17_req2[1], arbin16_req2[1], arbin15_req2[1], arbin14_req2[1],
    arbin13_req2[1], arbin12_req2[1], arbin11_req2[1], arbin10_req2[1],
    arbin09_req2[1], arbin08_req2[1], arbin07_req2[1], arbin06_req2[1],
    arbin05_req2[1], arbin04_req2[1], arbin03_req2[1], arbin02_req2[1],
    arbin01_req2[1], arbin00_req2[1]};

  assign arbout02_req2 = {
    arbin21_req2[2], arbin20_req2[2], arbin19_req2[2], arbin18_req2[2],
    arbin17_req2[2], arbin16_req2[2], arbin15_req2[2], arbin14_req2[2],
    arbin13_req2[2], arbin12_req2[2], arbin11_req2[2], arbin10_req2[2],
    arbin09_req2[2], arbin08_req2[2], arbin07_req2[2], arbin06_req2[2],
    arbin05_req2[2], arbin04_req2[2], arbin03_req2[2], arbin02_req2[2],
    arbin01_req2[2], arbin00_req2[2]};

  assign arbout03_req2 = {
    arbin21_req2[3], arbin20_req2[3], arbin19_req2[3], arbin18_req2[3],
    arbin17_req2[3], arbin16_req2[3], arbin15_req2[3], arbin14_req2[3],
    arbin13_req2[3], arbin12_req2[3], arbin11_req2[3], arbin10_req2[3],
    arbin09_req2[3], arbin08_req2[3], arbin07_req2[3], arbin06_req2[3],
    arbin05_req2[3], arbin04_req2[3], arbin03_req2[3], arbin02_req2[3],
    arbin01_req2[3], arbin00_req2[3]};

  assign arbout04_req2 = {
    arbin21_req2[4], arbin20_req2[4], arbin19_req2[4], arbin18_req2[4],
    arbin17_req2[4], arbin16_req2[4], arbin15_req2[4], arbin14_req2[4],
    arbin13_req2[4], arbin12_req2[4], arbin11_req2[4], arbin10_req2[4],
    arbin09_req2[4], arbin08_req2[4], arbin07_req2[4], arbin06_req2[4],
    arbin05_req2[4], arbin04_req2[4], arbin03_req2[4], arbin02_req2[4],
    arbin01_req2[4], arbin00_req2[4]};

  assign arbout05_req2 = {
    arbin21_req2[5], arbin20_req2[5], arbin19_req2[5], arbin18_req2[5],
    arbin17_req2[5], arbin16_req2[5], arbin15_req2[5], arbin14_req2[5],
    arbin13_req2[5], arbin12_req2[5], arbin11_req2[5], arbin10_req2[5],
    arbin09_req2[5], arbin08_req2[5], arbin07_req2[5], arbin06_req2[5],
    arbin05_req2[5], arbin04_req2[5], arbin03_req2[5], arbin02_req2[5],
    arbin01_req2[5], arbin00_req2[5]};

  assign arbout06_req2 = {
    arbin21_req2[6], arbin20_req2[6], arbin19_req2[6], arbin18_req2[6],
    arbin17_req2[6], arbin16_req2[6], arbin15_req2[6], arbin14_req2[6],
    arbin13_req2[6], arbin12_req2[6], arbin11_req2[6], arbin10_req2[6],
    arbin09_req2[6], arbin08_req2[6], arbin07_req2[6], arbin06_req2[6],
    arbin05_req2[6], arbin04_req2[6], arbin03_req2[6], arbin02_req2[6],
    arbin01_req2[6], arbin00_req2[6]};

  assign arbout07_req2 = {
    arbin21_req2[7], arbin20_req2[7], arbin19_req2[7], arbin18_req2[7],
    arbin17_req2[7], arbin16_req2[7], arbin15_req2[7], arbin14_req2[7],
    arbin13_req2[7], arbin12_req2[7], arbin11_req2[7], arbin10_req2[7],
    arbin09_req2[7], arbin08_req2[7], arbin07_req2[7], arbin06_req2[7],
    arbin05_req2[7], arbin04_req2[7], arbin03_req2[7], arbin02_req2[7],
    arbin01_req2[7], arbin00_req2[7]};

  assign arbout08_req2 = {
    arbin21_req2[8], arbin20_req2[8], arbin19_req2[8], arbin18_req2[8],
    arbin17_req2[8], arbin16_req2[8], arbin15_req2[8], arbin14_req2[8],
    arbin13_req2[8], arbin12_req2[8], arbin11_req2[8], arbin10_req2[8],
    arbin09_req2[8], arbin08_req2[8], arbin07_req2[8], arbin06_req2[8],
    arbin05_req2[8], arbin04_req2[8], arbin03_req2[8], arbin02_req2[8],
    arbin01_req2[8], arbin00_req2[8]};

  assign arbout09_req2 = {
    arbin21_req2[9], arbin20_req2[9], arbin19_req2[9], arbin18_req2[9],
    arbin17_req2[9], arbin16_req2[9], arbin15_req2[9], arbin14_req2[9],
    arbin13_req2[9], arbin12_req2[9], arbin11_req2[9], arbin10_req2[9],
    arbin09_req2[9], arbin08_req2[9], arbin07_req2[9], arbin06_req2[9],
    arbin05_req2[9], arbin04_req2[9], arbin03_req2[9], arbin02_req2[9],
    arbin01_req2[9], arbin00_req2[9]};

  assign arbout10_req2 = {
    arbin21_req2[10], arbin20_req2[10], arbin19_req2[10], arbin18_req2[10],
    arbin17_req2[10], arbin16_req2[10], arbin15_req2[10], arbin14_req2[10],
    arbin13_req2[10], arbin12_req2[10], arbin11_req2[10], arbin10_req2[10],
    arbin09_req2[10], arbin08_req2[10], arbin07_req2[10], arbin06_req2[10],
    arbin05_req2[10], arbin04_req2[10], arbin03_req2[10], arbin02_req2[10],
    arbin01_req2[10], arbin00_req2[10]};

  assign arbout11_req2 = {
    arbin21_req2[11], arbin20_req2[11], arbin19_req2[11], arbin18_req2[11],
    arbin17_req2[11], arbin16_req2[11], arbin15_req2[11], arbin14_req2[11],
    arbin13_req2[11], arbin12_req2[11], arbin11_req2[11], arbin10_req2[11],
    arbin09_req2[11], arbin08_req2[11], arbin07_req2[11], arbin06_req2[11],
    arbin05_req2[11], arbin04_req2[11], arbin03_req2[11], arbin02_req2[11],
    arbin01_req2[11], arbin00_req2[11]};

  assign arbout12_req2 = {
    arbin21_req2[12], arbin20_req2[12], arbin19_req2[12], arbin18_req2[12],
    arbin17_req2[12], arbin16_req2[12], arbin15_req2[12], arbin14_req2[12],
    arbin13_req2[12], arbin12_req2[12], arbin11_req2[12], arbin10_req2[12],
    arbin09_req2[12], arbin08_req2[12], arbin07_req2[12], arbin06_req2[12],
    arbin05_req2[12], arbin04_req2[12], arbin03_req2[12], arbin02_req2[12],
    arbin01_req2[12], arbin00_req2[12]};

  assign arbout13_req2 = {
    arbin21_req2[13], arbin20_req2[13], arbin19_req2[13], arbin18_req2[13],
    arbin17_req2[13], arbin16_req2[13], arbin15_req2[13], arbin14_req2[13],
    arbin13_req2[13], arbin12_req2[13], arbin11_req2[13], arbin10_req2[13],
    arbin09_req2[13], arbin08_req2[13], arbin07_req2[13], arbin06_req2[13],
    arbin05_req2[13], arbin04_req2[13], arbin03_req2[13], arbin02_req2[13],
    arbin01_req2[13], arbin00_req2[13]};

  assign arbout14_req2 = {
    arbin21_req2[14], arbin20_req2[14], arbin19_req2[14], arbin18_req2[14],
    arbin17_req2[14], arbin16_req2[14], arbin15_req2[14], arbin14_req2[14],
    arbin13_req2[14], arbin12_req2[14], arbin11_req2[14], arbin10_req2[14],
    arbin09_req2[14], arbin08_req2[14], arbin07_req2[14], arbin06_req2[14],
    arbin05_req2[14], arbin04_req2[14], arbin03_req2[14], arbin02_req2[14],
    arbin01_req2[14], arbin00_req2[14]};

  assign arbout15_req2 = {
    arbin21_req2[15], arbin20_req2[15], arbin19_req2[15], arbin18_req2[15],
    arbin17_req2[15], arbin16_req2[15], arbin15_req2[15], arbin14_req2[15],
    arbin13_req2[15], arbin12_req2[15], arbin11_req2[15], arbin10_req2[15],
    arbin09_req2[15], arbin08_req2[15], arbin07_req2[15], arbin06_req2[15],
    arbin05_req2[15], arbin04_req2[15], arbin03_req2[15], arbin02_req2[15],
    arbin01_req2[15], arbin00_req2[15]};

  assign arbout16_req2 = {
    arbin21_req2[16], arbin20_req2[16], arbin19_req2[16], arbin18_req2[16],
    arbin17_req2[16], arbin16_req2[16], arbin15_req2[16], arbin14_req2[16],
    arbin13_req2[16], arbin12_req2[16], arbin11_req2[16], arbin10_req2[16],
    arbin09_req2[16], arbin08_req2[16], arbin07_req2[16], arbin06_req2[16],
    arbin05_req2[16], arbin04_req2[16], arbin03_req2[16], arbin02_req2[16],
    arbin01_req2[16], arbin00_req2[16]};

  assign arbout17_req2 = {
    arbin21_req2[17], arbin20_req2[17], arbin19_req2[17], arbin18_req2[17],
    arbin17_req2[17], arbin16_req2[17], arbin15_req2[17], arbin14_req2[17],
    arbin13_req2[17], arbin12_req2[17], arbin11_req2[17], arbin10_req2[17],
    arbin09_req2[17], arbin08_req2[17], arbin07_req2[17], arbin06_req2[17],
    arbin05_req2[17], arbin04_req2[17], arbin03_req2[17], arbin02_req2[17],
    arbin01_req2[17], arbin00_req2[17]};

  assign arbout18_req2 = {
    arbin21_req2[18], arbin20_req2[18], arbin19_req2[18], arbin18_req2[18],
    arbin17_req2[18], arbin16_req2[18], arbin15_req2[18], arbin14_req2[18],
    arbin13_req2[18], arbin12_req2[18], arbin11_req2[18], arbin10_req2[18],
    arbin09_req2[18], arbin08_req2[18], arbin07_req2[18], arbin06_req2[18],
    arbin05_req2[18], arbin04_req2[18], arbin03_req2[18], arbin02_req2[18],
    arbin01_req2[18], arbin00_req2[18]};

  assign arbout19_req2 = {
    arbin21_req2[19], arbin20_req2[19], arbin19_req2[19], arbin18_req2[19],
    arbin17_req2[19], arbin16_req2[19], arbin15_req2[19], arbin14_req2[19],
    arbin13_req2[19], arbin12_req2[19], arbin11_req2[19], arbin10_req2[19],
    arbin09_req2[19], arbin08_req2[19], arbin07_req2[19], arbin06_req2[19],
    arbin05_req2[19], arbin04_req2[19], arbin03_req2[19], arbin02_req2[19],
    arbin01_req2[19], arbin00_req2[19]};

  assign arbout20_req2 = {
    arbin21_req2[20], arbin20_req2[20], arbin19_req2[20], arbin18_req2[20],
    arbin17_req2[20], arbin16_req2[20], arbin15_req2[20], arbin14_req2[20],
    arbin13_req2[20], arbin12_req2[20], arbin11_req2[20], arbin10_req2[20],
    arbin09_req2[20], arbin08_req2[20], arbin07_req2[20], arbin06_req2[20],
    arbin05_req2[20], arbin04_req2[20], arbin03_req2[20], arbin02_req2[20],
    arbin01_req2[20], arbin00_req2[20]};

  assign arbout21_req2 = {
    arbin21_req2[21], arbin20_req2[21], arbin19_req2[21], arbin18_req2[21],
    arbin17_req2[21], arbin16_req2[21], arbin15_req2[21], arbin14_req2[21],
    arbin13_req2[21], arbin12_req2[21], arbin11_req2[21], arbin10_req2[21],
    arbin09_req2[21], arbin08_req2[21], arbin07_req2[21], arbin06_req2[21],
    arbin05_req2[21], arbin04_req2[21], arbin03_req2[21], arbin02_req2[21],
    arbin01_req2[21], arbin00_req2[21]};

  
  // ==========================================================================
  // Grant stiching
  // ==========================================================================
  assign arbin00_gnt0 = {
    arbout21_gnt0[0], arbout20_gnt0[0], arbout19_gnt0[0], arbout18_gnt0[0],
    arbout17_gnt0[0], arbout16_gnt0[0], arbout15_gnt0[0], arbout14_gnt0[0],
    arbout13_gnt0[0], arbout12_gnt0[0], arbout11_gnt0[0], arbout10_gnt0[0],
    arbout09_gnt0[0], arbout08_gnt0[0], arbout07_gnt0[0], arbout06_gnt0[0],
    arbout05_gnt0[0], arbout04_gnt0[0], arbout03_gnt0[0], arbout02_gnt0[0],
    arbout01_gnt0[0], arbout00_gnt0[0]};

  assign arbin01_gnt0 = {
    arbout21_gnt0[1], arbout20_gnt0[1], arbout19_gnt0[1], arbout18_gnt0[1],
    arbout17_gnt0[1], arbout16_gnt0[1], arbout15_gnt0[1], arbout14_gnt0[1],
    arbout13_gnt0[1], arbout12_gnt0[1], arbout11_gnt0[1], arbout10_gnt0[1],
    arbout09_gnt0[1], arbout08_gnt0[1], arbout07_gnt0[1], arbout06_gnt0[1],
    arbout05_gnt0[1], arbout04_gnt0[1], arbout03_gnt0[1], arbout02_gnt0[1],
    arbout01_gnt0[1], arbout00_gnt0[1]};

  assign arbin02_gnt0 = {
    arbout21_gnt0[2], arbout20_gnt0[2], arbout19_gnt0[2], arbout18_gnt0[2],
    arbout17_gnt0[2], arbout16_gnt0[2], arbout15_gnt0[2], arbout14_gnt0[2],
    arbout13_gnt0[2], arbout12_gnt0[2], arbout11_gnt0[2], arbout10_gnt0[2],
    arbout09_gnt0[2], arbout08_gnt0[2], arbout07_gnt0[2], arbout06_gnt0[2],
    arbout05_gnt0[2], arbout04_gnt0[2], arbout03_gnt0[2], arbout02_gnt0[2],
    arbout01_gnt0[2], arbout00_gnt0[2]};

  assign arbin03_gnt0 = {
    arbout21_gnt0[3], arbout20_gnt0[3], arbout19_gnt0[3], arbout18_gnt0[3],
    arbout17_gnt0[3], arbout16_gnt0[3], arbout15_gnt0[3], arbout14_gnt0[3],
    arbout13_gnt0[3], arbout12_gnt0[3], arbout11_gnt0[3], arbout10_gnt0[3],
    arbout09_gnt0[3], arbout08_gnt0[3], arbout07_gnt0[3], arbout06_gnt0[3],
    arbout05_gnt0[3], arbout04_gnt0[3], arbout03_gnt0[3], arbout02_gnt0[3],
    arbout01_gnt0[3], arbout00_gnt0[3]};

  assign arbin04_gnt0 = {
    arbout21_gnt0[4], arbout20_gnt0[4], arbout19_gnt0[4], arbout18_gnt0[4],
    arbout17_gnt0[4], arbout16_gnt0[4], arbout15_gnt0[4], arbout14_gnt0[4],
    arbout13_gnt0[4], arbout12_gnt0[4], arbout11_gnt0[4], arbout10_gnt0[4],
    arbout09_gnt0[4], arbout08_gnt0[4], arbout07_gnt0[4], arbout06_gnt0[4],
    arbout05_gnt0[4], arbout04_gnt0[4], arbout03_gnt0[4], arbout02_gnt0[4],
    arbout01_gnt0[4], arbout00_gnt0[4]};

  assign arbin05_gnt0 = {
    arbout21_gnt0[5], arbout20_gnt0[5], arbout19_gnt0[5], arbout18_gnt0[5],
    arbout17_gnt0[5], arbout16_gnt0[5], arbout15_gnt0[5], arbout14_gnt0[5],
    arbout13_gnt0[5], arbout12_gnt0[5], arbout11_gnt0[5], arbout10_gnt0[5],
    arbout09_gnt0[5], arbout08_gnt0[5], arbout07_gnt0[5], arbout06_gnt0[5],
    arbout05_gnt0[5], arbout04_gnt0[5], arbout03_gnt0[5], arbout02_gnt0[5],
    arbout01_gnt0[5], arbout00_gnt0[5]};

  assign arbin06_gnt0 = {
    arbout21_gnt0[6], arbout20_gnt0[6], arbout19_gnt0[6], arbout18_gnt0[6],
    arbout17_gnt0[6], arbout16_gnt0[6], arbout15_gnt0[6], arbout14_gnt0[6],
    arbout13_gnt0[6], arbout12_gnt0[6], arbout11_gnt0[6], arbout10_gnt0[6],
    arbout09_gnt0[6], arbout08_gnt0[6], arbout07_gnt0[6], arbout06_gnt0[6],
    arbout05_gnt0[6], arbout04_gnt0[6], arbout03_gnt0[6], arbout02_gnt0[6],
    arbout01_gnt0[6], arbout00_gnt0[6]};

  assign arbin07_gnt0 = {
    arbout21_gnt0[7], arbout20_gnt0[7], arbout19_gnt0[7], arbout18_gnt0[7],
    arbout17_gnt0[7], arbout16_gnt0[7], arbout15_gnt0[7], arbout14_gnt0[7],
    arbout13_gnt0[7], arbout12_gnt0[7], arbout11_gnt0[7], arbout10_gnt0[7],
    arbout09_gnt0[7], arbout08_gnt0[7], arbout07_gnt0[7], arbout06_gnt0[7],
    arbout05_gnt0[7], arbout04_gnt0[7], arbout03_gnt0[7], arbout02_gnt0[7],
    arbout01_gnt0[7], arbout00_gnt0[7]};

  assign arbin08_gnt0 = {
    arbout21_gnt0[8], arbout20_gnt0[8], arbout19_gnt0[8], arbout18_gnt0[8],
    arbout17_gnt0[8], arbout16_gnt0[8], arbout15_gnt0[8], arbout14_gnt0[8],
    arbout13_gnt0[8], arbout12_gnt0[8], arbout11_gnt0[8], arbout10_gnt0[8],
    arbout09_gnt0[8], arbout08_gnt0[8], arbout07_gnt0[8], arbout06_gnt0[8],
    arbout05_gnt0[8], arbout04_gnt0[8], arbout03_gnt0[8], arbout02_gnt0[8],
    arbout01_gnt0[8], arbout00_gnt0[8]};

  assign arbin09_gnt0 = {
    arbout21_gnt0[9], arbout20_gnt0[9], arbout19_gnt0[9], arbout18_gnt0[9],
    arbout17_gnt0[9], arbout16_gnt0[9], arbout15_gnt0[9], arbout14_gnt0[9],
    arbout13_gnt0[9], arbout12_gnt0[9], arbout11_gnt0[9], arbout10_gnt0[9],
    arbout09_gnt0[9], arbout08_gnt0[9], arbout07_gnt0[9], arbout06_gnt0[9],
    arbout05_gnt0[9], arbout04_gnt0[9], arbout03_gnt0[9], arbout02_gnt0[9],
    arbout01_gnt0[9], arbout00_gnt0[9]};

  assign arbin10_gnt0 = {
    arbout21_gnt0[10], arbout20_gnt0[10], arbout19_gnt0[10], arbout18_gnt0[10],
    arbout17_gnt0[10], arbout16_gnt0[10], arbout15_gnt0[10], arbout14_gnt0[10],
    arbout13_gnt0[10], arbout12_gnt0[10], arbout11_gnt0[10], arbout10_gnt0[10],
    arbout09_gnt0[10], arbout08_gnt0[10], arbout07_gnt0[10], arbout06_gnt0[10],
    arbout05_gnt0[10], arbout04_gnt0[10], arbout03_gnt0[10], arbout02_gnt0[10],
    arbout01_gnt0[10], arbout00_gnt0[10]};

  assign arbin11_gnt0 = {
    arbout21_gnt0[11], arbout20_gnt0[11], arbout19_gnt0[11], arbout18_gnt0[11],
    arbout17_gnt0[11], arbout16_gnt0[11], arbout15_gnt0[11], arbout14_gnt0[11],
    arbout13_gnt0[11], arbout12_gnt0[11], arbout11_gnt0[11], arbout10_gnt0[11],
    arbout09_gnt0[11], arbout08_gnt0[11], arbout07_gnt0[11], arbout06_gnt0[11],
    arbout05_gnt0[11], arbout04_gnt0[11], arbout03_gnt0[11], arbout02_gnt0[11],
    arbout01_gnt0[11], arbout00_gnt0[11]};

  assign arbin12_gnt0 = {
    arbout21_gnt0[12], arbout20_gnt0[12], arbout19_gnt0[12], arbout18_gnt0[12],
    arbout17_gnt0[12], arbout16_gnt0[12], arbout15_gnt0[12], arbout14_gnt0[12],
    arbout13_gnt0[12], arbout12_gnt0[12], arbout11_gnt0[12], arbout10_gnt0[12],
    arbout09_gnt0[12], arbout08_gnt0[12], arbout07_gnt0[12], arbout06_gnt0[12],
    arbout05_gnt0[12], arbout04_gnt0[12], arbout03_gnt0[12], arbout02_gnt0[12],
    arbout01_gnt0[12], arbout00_gnt0[12]};

  assign arbin13_gnt0 = {
    arbout21_gnt0[13], arbout20_gnt0[13], arbout19_gnt0[13], arbout18_gnt0[13],
    arbout17_gnt0[13], arbout16_gnt0[13], arbout15_gnt0[13], arbout14_gnt0[13],
    arbout13_gnt0[13], arbout12_gnt0[13], arbout11_gnt0[13], arbout10_gnt0[13],
    arbout09_gnt0[13], arbout08_gnt0[13], arbout07_gnt0[13], arbout06_gnt0[13],
    arbout05_gnt0[13], arbout04_gnt0[13], arbout03_gnt0[13], arbout02_gnt0[13],
    arbout01_gnt0[13], arbout00_gnt0[13]};

  assign arbin14_gnt0 = {
    arbout21_gnt0[14], arbout20_gnt0[14], arbout19_gnt0[14], arbout18_gnt0[14],
    arbout17_gnt0[14], arbout16_gnt0[14], arbout15_gnt0[14], arbout14_gnt0[14],
    arbout13_gnt0[14], arbout12_gnt0[14], arbout11_gnt0[14], arbout10_gnt0[14],
    arbout09_gnt0[14], arbout08_gnt0[14], arbout07_gnt0[14], arbout06_gnt0[14],
    arbout05_gnt0[14], arbout04_gnt0[14], arbout03_gnt0[14], arbout02_gnt0[14],
    arbout01_gnt0[14], arbout00_gnt0[14]};

  assign arbin15_gnt0 = {
    arbout21_gnt0[15], arbout20_gnt0[15], arbout19_gnt0[15], arbout18_gnt0[15],
    arbout17_gnt0[15], arbout16_gnt0[15], arbout15_gnt0[15], arbout14_gnt0[15],
    arbout13_gnt0[15], arbout12_gnt0[15], arbout11_gnt0[15], arbout10_gnt0[15],
    arbout09_gnt0[15], arbout08_gnt0[15], arbout07_gnt0[15], arbout06_gnt0[15],
    arbout05_gnt0[15], arbout04_gnt0[15], arbout03_gnt0[15], arbout02_gnt0[15],
    arbout01_gnt0[15], arbout00_gnt0[15]};

  assign arbin16_gnt0 = {
    arbout21_gnt0[16], arbout20_gnt0[16], arbout19_gnt0[16], arbout18_gnt0[16],
    arbout17_gnt0[16], arbout16_gnt0[16], arbout15_gnt0[16], arbout14_gnt0[16],
    arbout13_gnt0[16], arbout12_gnt0[16], arbout11_gnt0[16], arbout10_gnt0[16],
    arbout09_gnt0[16], arbout08_gnt0[16], arbout07_gnt0[16], arbout06_gnt0[16],
    arbout05_gnt0[16], arbout04_gnt0[16], arbout03_gnt0[16], arbout02_gnt0[16],
    arbout01_gnt0[16], arbout00_gnt0[16]};

  assign arbin17_gnt0 = {
    arbout21_gnt0[17], arbout20_gnt0[17], arbout19_gnt0[17], arbout18_gnt0[17],
    arbout17_gnt0[17], arbout16_gnt0[17], arbout15_gnt0[17], arbout14_gnt0[17],
    arbout13_gnt0[17], arbout12_gnt0[17], arbout11_gnt0[17], arbout10_gnt0[17],
    arbout09_gnt0[17], arbout08_gnt0[17], arbout07_gnt0[17], arbout06_gnt0[17],
    arbout05_gnt0[17], arbout04_gnt0[17], arbout03_gnt0[17], arbout02_gnt0[17],
    arbout01_gnt0[17], arbout00_gnt0[17]};

  assign arbin18_gnt0 = {
    arbout21_gnt0[18], arbout20_gnt0[18], arbout19_gnt0[18], arbout18_gnt0[18],
    arbout17_gnt0[18], arbout16_gnt0[18], arbout15_gnt0[18], arbout14_gnt0[18],
    arbout13_gnt0[18], arbout12_gnt0[18], arbout11_gnt0[18], arbout10_gnt0[18],
    arbout09_gnt0[18], arbout08_gnt0[18], arbout07_gnt0[18], arbout06_gnt0[18],
    arbout05_gnt0[18], arbout04_gnt0[18], arbout03_gnt0[18], arbout02_gnt0[18],
    arbout01_gnt0[18], arbout00_gnt0[18]};

  assign arbin19_gnt0 = {
    arbout21_gnt0[19], arbout20_gnt0[19], arbout19_gnt0[19], arbout18_gnt0[19],
    arbout17_gnt0[19], arbout16_gnt0[19], arbout15_gnt0[19], arbout14_gnt0[19],
    arbout13_gnt0[19], arbout12_gnt0[19], arbout11_gnt0[19], arbout10_gnt0[19],
    arbout09_gnt0[19], arbout08_gnt0[19], arbout07_gnt0[19], arbout06_gnt0[19],
    arbout05_gnt0[19], arbout04_gnt0[19], arbout03_gnt0[19], arbout02_gnt0[19],
    arbout01_gnt0[19], arbout00_gnt0[19]};

  assign arbin20_gnt0 = {
    arbout21_gnt0[20], arbout20_gnt0[20], arbout19_gnt0[20], arbout18_gnt0[20],
    arbout17_gnt0[20], arbout16_gnt0[20], arbout15_gnt0[20], arbout14_gnt0[20],
    arbout13_gnt0[20], arbout12_gnt0[20], arbout11_gnt0[20], arbout10_gnt0[20],
    arbout09_gnt0[20], arbout08_gnt0[20], arbout07_gnt0[20], arbout06_gnt0[20],
    arbout05_gnt0[20], arbout04_gnt0[20], arbout03_gnt0[20], arbout02_gnt0[20],
    arbout01_gnt0[20], arbout00_gnt0[20]};

  assign arbin21_gnt0 = {
    arbout21_gnt0[21], arbout20_gnt0[21], arbout19_gnt0[21], arbout18_gnt0[21],
    arbout17_gnt0[21], arbout16_gnt0[21], arbout15_gnt0[21], arbout14_gnt0[21],
    arbout13_gnt0[21], arbout12_gnt0[21], arbout11_gnt0[21], arbout10_gnt0[21],
    arbout09_gnt0[21], arbout08_gnt0[21], arbout07_gnt0[21], arbout06_gnt0[21],
    arbout05_gnt0[21], arbout04_gnt0[21], arbout03_gnt0[21], arbout02_gnt0[21],
    arbout01_gnt0[21], arbout00_gnt0[21]};

  assign arbin00_gnt1 = {
    arbout21_gnt1[0], arbout20_gnt1[0], arbout19_gnt1[0], arbout18_gnt1[0],
    arbout17_gnt1[0], arbout16_gnt1[0], arbout15_gnt1[0], arbout14_gnt1[0],
    arbout13_gnt1[0], arbout12_gnt1[0], arbout11_gnt1[0], arbout10_gnt1[0],
    arbout09_gnt1[0], arbout08_gnt1[0], arbout07_gnt1[0], arbout06_gnt1[0],
    arbout05_gnt1[0], arbout04_gnt1[0], arbout03_gnt1[0], arbout02_gnt1[0],
    arbout01_gnt1[0], arbout00_gnt1[0]};

  assign arbin01_gnt1 = {
    arbout21_gnt1[1], arbout20_gnt1[1], arbout19_gnt1[1], arbout18_gnt1[1],
    arbout17_gnt1[1], arbout16_gnt1[1], arbout15_gnt1[1], arbout14_gnt1[1],
    arbout13_gnt1[1], arbout12_gnt1[1], arbout11_gnt1[1], arbout10_gnt1[1],
    arbout09_gnt1[1], arbout08_gnt1[1], arbout07_gnt1[1], arbout06_gnt1[1],
    arbout05_gnt1[1], arbout04_gnt1[1], arbout03_gnt1[1], arbout02_gnt1[1],
    arbout01_gnt1[1], arbout00_gnt1[1]};

  assign arbin02_gnt1 = {
    arbout21_gnt1[2], arbout20_gnt1[2], arbout19_gnt1[2], arbout18_gnt1[2],
    arbout17_gnt1[2], arbout16_gnt1[2], arbout15_gnt1[2], arbout14_gnt1[2],
    arbout13_gnt1[2], arbout12_gnt1[2], arbout11_gnt1[2], arbout10_gnt1[2],
    arbout09_gnt1[2], arbout08_gnt1[2], arbout07_gnt1[2], arbout06_gnt1[2],
    arbout05_gnt1[2], arbout04_gnt1[2], arbout03_gnt1[2], arbout02_gnt1[2],
    arbout01_gnt1[2], arbout00_gnt1[2]};

  assign arbin03_gnt1 = {
    arbout21_gnt1[3], arbout20_gnt1[3], arbout19_gnt1[3], arbout18_gnt1[3],
    arbout17_gnt1[3], arbout16_gnt1[3], arbout15_gnt1[3], arbout14_gnt1[3],
    arbout13_gnt1[3], arbout12_gnt1[3], arbout11_gnt1[3], arbout10_gnt1[3],
    arbout09_gnt1[3], arbout08_gnt1[3], arbout07_gnt1[3], arbout06_gnt1[3],
    arbout05_gnt1[3], arbout04_gnt1[3], arbout03_gnt1[3], arbout02_gnt1[3],
    arbout01_gnt1[3], arbout00_gnt1[3]};

  assign arbin04_gnt1 = {
    arbout21_gnt1[4], arbout20_gnt1[4], arbout19_gnt1[4], arbout18_gnt1[4],
    arbout17_gnt1[4], arbout16_gnt1[4], arbout15_gnt1[4], arbout14_gnt1[4],
    arbout13_gnt1[4], arbout12_gnt1[4], arbout11_gnt1[4], arbout10_gnt1[4],
    arbout09_gnt1[4], arbout08_gnt1[4], arbout07_gnt1[4], arbout06_gnt1[4],
    arbout05_gnt1[4], arbout04_gnt1[4], arbout03_gnt1[4], arbout02_gnt1[4],
    arbout01_gnt1[4], arbout00_gnt1[4]};

  assign arbin05_gnt1 = {
    arbout21_gnt1[5], arbout20_gnt1[5], arbout19_gnt1[5], arbout18_gnt1[5],
    arbout17_gnt1[5], arbout16_gnt1[5], arbout15_gnt1[5], arbout14_gnt1[5],
    arbout13_gnt1[5], arbout12_gnt1[5], arbout11_gnt1[5], arbout10_gnt1[5],
    arbout09_gnt1[5], arbout08_gnt1[5], arbout07_gnt1[5], arbout06_gnt1[5],
    arbout05_gnt1[5], arbout04_gnt1[5], arbout03_gnt1[5], arbout02_gnt1[5],
    arbout01_gnt1[5], arbout00_gnt1[5]};

  assign arbin06_gnt1 = {
    arbout21_gnt1[6], arbout20_gnt1[6], arbout19_gnt1[6], arbout18_gnt1[6],
    arbout17_gnt1[6], arbout16_gnt1[6], arbout15_gnt1[6], arbout14_gnt1[6],
    arbout13_gnt1[6], arbout12_gnt1[6], arbout11_gnt1[6], arbout10_gnt1[6],
    arbout09_gnt1[6], arbout08_gnt1[6], arbout07_gnt1[6], arbout06_gnt1[6],
    arbout05_gnt1[6], arbout04_gnt1[6], arbout03_gnt1[6], arbout02_gnt1[6],
    arbout01_gnt1[6], arbout00_gnt1[6]};

  assign arbin07_gnt1 = {
    arbout21_gnt1[7], arbout20_gnt1[7], arbout19_gnt1[7], arbout18_gnt1[7],
    arbout17_gnt1[7], arbout16_gnt1[7], arbout15_gnt1[7], arbout14_gnt1[7],
    arbout13_gnt1[7], arbout12_gnt1[7], arbout11_gnt1[7], arbout10_gnt1[7],
    arbout09_gnt1[7], arbout08_gnt1[7], arbout07_gnt1[7], arbout06_gnt1[7],
    arbout05_gnt1[7], arbout04_gnt1[7], arbout03_gnt1[7], arbout02_gnt1[7],
    arbout01_gnt1[7], arbout00_gnt1[7]};

  assign arbin08_gnt1 = {
    arbout21_gnt1[8], arbout20_gnt1[8], arbout19_gnt1[8], arbout18_gnt1[8],
    arbout17_gnt1[8], arbout16_gnt1[8], arbout15_gnt1[8], arbout14_gnt1[8],
    arbout13_gnt1[8], arbout12_gnt1[8], arbout11_gnt1[8], arbout10_gnt1[8],
    arbout09_gnt1[8], arbout08_gnt1[8], arbout07_gnt1[8], arbout06_gnt1[8],
    arbout05_gnt1[8], arbout04_gnt1[8], arbout03_gnt1[8], arbout02_gnt1[8],
    arbout01_gnt1[8], arbout00_gnt1[8]};

  assign arbin09_gnt1 = {
    arbout21_gnt1[9], arbout20_gnt1[9], arbout19_gnt1[9], arbout18_gnt1[9],
    arbout17_gnt1[9], arbout16_gnt1[9], arbout15_gnt1[9], arbout14_gnt1[9],
    arbout13_gnt1[9], arbout12_gnt1[9], arbout11_gnt1[9], arbout10_gnt1[9],
    arbout09_gnt1[9], arbout08_gnt1[9], arbout07_gnt1[9], arbout06_gnt1[9],
    arbout05_gnt1[9], arbout04_gnt1[9], arbout03_gnt1[9], arbout02_gnt1[9],
    arbout01_gnt1[9], arbout00_gnt1[9]};

  assign arbin10_gnt1 = {
    arbout21_gnt1[10], arbout20_gnt1[10], arbout19_gnt1[10], arbout18_gnt1[10],
    arbout17_gnt1[10], arbout16_gnt1[10], arbout15_gnt1[10], arbout14_gnt1[10],
    arbout13_gnt1[10], arbout12_gnt1[10], arbout11_gnt1[10], arbout10_gnt1[10],
    arbout09_gnt1[10], arbout08_gnt1[10], arbout07_gnt1[10], arbout06_gnt1[10],
    arbout05_gnt1[10], arbout04_gnt1[10], arbout03_gnt1[10], arbout02_gnt1[10],
    arbout01_gnt1[10], arbout00_gnt1[10]};

  assign arbin11_gnt1 = {
    arbout21_gnt1[11], arbout20_gnt1[11], arbout19_gnt1[11], arbout18_gnt1[11],
    arbout17_gnt1[11], arbout16_gnt1[11], arbout15_gnt1[11], arbout14_gnt1[11],
    arbout13_gnt1[11], arbout12_gnt1[11], arbout11_gnt1[11], arbout10_gnt1[11],
    arbout09_gnt1[11], arbout08_gnt1[11], arbout07_gnt1[11], arbout06_gnt1[11],
    arbout05_gnt1[11], arbout04_gnt1[11], arbout03_gnt1[11], arbout02_gnt1[11],
    arbout01_gnt1[11], arbout00_gnt1[11]};

  assign arbin12_gnt1 = {
    arbout21_gnt1[12], arbout20_gnt1[12], arbout19_gnt1[12], arbout18_gnt1[12],
    arbout17_gnt1[12], arbout16_gnt1[12], arbout15_gnt1[12], arbout14_gnt1[12],
    arbout13_gnt1[12], arbout12_gnt1[12], arbout11_gnt1[12], arbout10_gnt1[12],
    arbout09_gnt1[12], arbout08_gnt1[12], arbout07_gnt1[12], arbout06_gnt1[12],
    arbout05_gnt1[12], arbout04_gnt1[12], arbout03_gnt1[12], arbout02_gnt1[12],
    arbout01_gnt1[12], arbout00_gnt1[12]};

  assign arbin13_gnt1 = {
    arbout21_gnt1[13], arbout20_gnt1[13], arbout19_gnt1[13], arbout18_gnt1[13],
    arbout17_gnt1[13], arbout16_gnt1[13], arbout15_gnt1[13], arbout14_gnt1[13],
    arbout13_gnt1[13], arbout12_gnt1[13], arbout11_gnt1[13], arbout10_gnt1[13],
    arbout09_gnt1[13], arbout08_gnt1[13], arbout07_gnt1[13], arbout06_gnt1[13],
    arbout05_gnt1[13], arbout04_gnt1[13], arbout03_gnt1[13], arbout02_gnt1[13],
    arbout01_gnt1[13], arbout00_gnt1[13]};

  assign arbin14_gnt1 = {
    arbout21_gnt1[14], arbout20_gnt1[14], arbout19_gnt1[14], arbout18_gnt1[14],
    arbout17_gnt1[14], arbout16_gnt1[14], arbout15_gnt1[14], arbout14_gnt1[14],
    arbout13_gnt1[14], arbout12_gnt1[14], arbout11_gnt1[14], arbout10_gnt1[14],
    arbout09_gnt1[14], arbout08_gnt1[14], arbout07_gnt1[14], arbout06_gnt1[14],
    arbout05_gnt1[14], arbout04_gnt1[14], arbout03_gnt1[14], arbout02_gnt1[14],
    arbout01_gnt1[14], arbout00_gnt1[14]};

  assign arbin15_gnt1 = {
    arbout21_gnt1[15], arbout20_gnt1[15], arbout19_gnt1[15], arbout18_gnt1[15],
    arbout17_gnt1[15], arbout16_gnt1[15], arbout15_gnt1[15], arbout14_gnt1[15],
    arbout13_gnt1[15], arbout12_gnt1[15], arbout11_gnt1[15], arbout10_gnt1[15],
    arbout09_gnt1[15], arbout08_gnt1[15], arbout07_gnt1[15], arbout06_gnt1[15],
    arbout05_gnt1[15], arbout04_gnt1[15], arbout03_gnt1[15], arbout02_gnt1[15],
    arbout01_gnt1[15], arbout00_gnt1[15]};

  assign arbin16_gnt1 = {
    arbout21_gnt1[16], arbout20_gnt1[16], arbout19_gnt1[16], arbout18_gnt1[16],
    arbout17_gnt1[16], arbout16_gnt1[16], arbout15_gnt1[16], arbout14_gnt1[16],
    arbout13_gnt1[16], arbout12_gnt1[16], arbout11_gnt1[16], arbout10_gnt1[16],
    arbout09_gnt1[16], arbout08_gnt1[16], arbout07_gnt1[16], arbout06_gnt1[16],
    arbout05_gnt1[16], arbout04_gnt1[16], arbout03_gnt1[16], arbout02_gnt1[16],
    arbout01_gnt1[16], arbout00_gnt1[16]};

  assign arbin17_gnt1 = {
    arbout21_gnt1[17], arbout20_gnt1[17], arbout19_gnt1[17], arbout18_gnt1[17],
    arbout17_gnt1[17], arbout16_gnt1[17], arbout15_gnt1[17], arbout14_gnt1[17],
    arbout13_gnt1[17], arbout12_gnt1[17], arbout11_gnt1[17], arbout10_gnt1[17],
    arbout09_gnt1[17], arbout08_gnt1[17], arbout07_gnt1[17], arbout06_gnt1[17],
    arbout05_gnt1[17], arbout04_gnt1[17], arbout03_gnt1[17], arbout02_gnt1[17],
    arbout01_gnt1[17], arbout00_gnt1[17]};

  assign arbin18_gnt1 = {
    arbout21_gnt1[18], arbout20_gnt1[18], arbout19_gnt1[18], arbout18_gnt1[18],
    arbout17_gnt1[18], arbout16_gnt1[18], arbout15_gnt1[18], arbout14_gnt1[18],
    arbout13_gnt1[18], arbout12_gnt1[18], arbout11_gnt1[18], arbout10_gnt1[18],
    arbout09_gnt1[18], arbout08_gnt1[18], arbout07_gnt1[18], arbout06_gnt1[18],
    arbout05_gnt1[18], arbout04_gnt1[18], arbout03_gnt1[18], arbout02_gnt1[18],
    arbout01_gnt1[18], arbout00_gnt1[18]};

  assign arbin19_gnt1 = {
    arbout21_gnt1[19], arbout20_gnt1[19], arbout19_gnt1[19], arbout18_gnt1[19],
    arbout17_gnt1[19], arbout16_gnt1[19], arbout15_gnt1[19], arbout14_gnt1[19],
    arbout13_gnt1[19], arbout12_gnt1[19], arbout11_gnt1[19], arbout10_gnt1[19],
    arbout09_gnt1[19], arbout08_gnt1[19], arbout07_gnt1[19], arbout06_gnt1[19],
    arbout05_gnt1[19], arbout04_gnt1[19], arbout03_gnt1[19], arbout02_gnt1[19],
    arbout01_gnt1[19], arbout00_gnt1[19]};

  assign arbin20_gnt1 = {
    arbout21_gnt1[20], arbout20_gnt1[20], arbout19_gnt1[20], arbout18_gnt1[20],
    arbout17_gnt1[20], arbout16_gnt1[20], arbout15_gnt1[20], arbout14_gnt1[20],
    arbout13_gnt1[20], arbout12_gnt1[20], arbout11_gnt1[20], arbout10_gnt1[20],
    arbout09_gnt1[20], arbout08_gnt1[20], arbout07_gnt1[20], arbout06_gnt1[20],
    arbout05_gnt1[20], arbout04_gnt1[20], arbout03_gnt1[20], arbout02_gnt1[20],
    arbout01_gnt1[20], arbout00_gnt1[20]};

  assign arbin21_gnt1 = {
    arbout21_gnt1[21], arbout20_gnt1[21], arbout19_gnt1[21], arbout18_gnt1[21],
    arbout17_gnt1[21], arbout16_gnt1[21], arbout15_gnt1[21], arbout14_gnt1[21],
    arbout13_gnt1[21], arbout12_gnt1[21], arbout11_gnt1[21], arbout10_gnt1[21],
    arbout09_gnt1[21], arbout08_gnt1[21], arbout07_gnt1[21], arbout06_gnt1[21],
    arbout05_gnt1[21], arbout04_gnt1[21], arbout03_gnt1[21], arbout02_gnt1[21],
    arbout01_gnt1[21], arbout00_gnt1[21]};

  assign arbin00_gnt2 = {
    arbout21_gnt2[0], arbout20_gnt2[0], arbout19_gnt2[0], arbout18_gnt2[0],
    arbout17_gnt2[0], arbout16_gnt2[0], arbout15_gnt2[0], arbout14_gnt2[0],
    arbout13_gnt2[0], arbout12_gnt2[0], arbout11_gnt2[0], arbout10_gnt2[0],
    arbout09_gnt2[0], arbout08_gnt2[0], arbout07_gnt2[0], arbout06_gnt2[0],
    arbout05_gnt2[0], arbout04_gnt2[0], arbout03_gnt2[0], arbout02_gnt2[0],
    arbout01_gnt2[0], arbout00_gnt2[0]};

  assign arbin01_gnt2 = {
    arbout21_gnt2[1], arbout20_gnt2[1], arbout19_gnt2[1], arbout18_gnt2[1],
    arbout17_gnt2[1], arbout16_gnt2[1], arbout15_gnt2[1], arbout14_gnt2[1],
    arbout13_gnt2[1], arbout12_gnt2[1], arbout11_gnt2[1], arbout10_gnt2[1],
    arbout09_gnt2[1], arbout08_gnt2[1], arbout07_gnt2[1], arbout06_gnt2[1],
    arbout05_gnt2[1], arbout04_gnt2[1], arbout03_gnt2[1], arbout02_gnt2[1],
    arbout01_gnt2[1], arbout00_gnt2[1]};

  assign arbin02_gnt2 = {
    arbout21_gnt2[2], arbout20_gnt2[2], arbout19_gnt2[2], arbout18_gnt2[2],
    arbout17_gnt2[2], arbout16_gnt2[2], arbout15_gnt2[2], arbout14_gnt2[2],
    arbout13_gnt2[2], arbout12_gnt2[2], arbout11_gnt2[2], arbout10_gnt2[2],
    arbout09_gnt2[2], arbout08_gnt2[2], arbout07_gnt2[2], arbout06_gnt2[2],
    arbout05_gnt2[2], arbout04_gnt2[2], arbout03_gnt2[2], arbout02_gnt2[2],
    arbout01_gnt2[2], arbout00_gnt2[2]};

  assign arbin03_gnt2 = {
    arbout21_gnt2[3], arbout20_gnt2[3], arbout19_gnt2[3], arbout18_gnt2[3],
    arbout17_gnt2[3], arbout16_gnt2[3], arbout15_gnt2[3], arbout14_gnt2[3],
    arbout13_gnt2[3], arbout12_gnt2[3], arbout11_gnt2[3], arbout10_gnt2[3],
    arbout09_gnt2[3], arbout08_gnt2[3], arbout07_gnt2[3], arbout06_gnt2[3],
    arbout05_gnt2[3], arbout04_gnt2[3], arbout03_gnt2[3], arbout02_gnt2[3],
    arbout01_gnt2[3], arbout00_gnt2[3]};

  assign arbin04_gnt2 = {
    arbout21_gnt2[4], arbout20_gnt2[4], arbout19_gnt2[4], arbout18_gnt2[4],
    arbout17_gnt2[4], arbout16_gnt2[4], arbout15_gnt2[4], arbout14_gnt2[4],
    arbout13_gnt2[4], arbout12_gnt2[4], arbout11_gnt2[4], arbout10_gnt2[4],
    arbout09_gnt2[4], arbout08_gnt2[4], arbout07_gnt2[4], arbout06_gnt2[4],
    arbout05_gnt2[4], arbout04_gnt2[4], arbout03_gnt2[4], arbout02_gnt2[4],
    arbout01_gnt2[4], arbout00_gnt2[4]};

  assign arbin05_gnt2 = {
    arbout21_gnt2[5], arbout20_gnt2[5], arbout19_gnt2[5], arbout18_gnt2[5],
    arbout17_gnt2[5], arbout16_gnt2[5], arbout15_gnt2[5], arbout14_gnt2[5],
    arbout13_gnt2[5], arbout12_gnt2[5], arbout11_gnt2[5], arbout10_gnt2[5],
    arbout09_gnt2[5], arbout08_gnt2[5], arbout07_gnt2[5], arbout06_gnt2[5],
    arbout05_gnt2[5], arbout04_gnt2[5], arbout03_gnt2[5], arbout02_gnt2[5],
    arbout01_gnt2[5], arbout00_gnt2[5]};

  assign arbin06_gnt2 = {
    arbout21_gnt2[6], arbout20_gnt2[6], arbout19_gnt2[6], arbout18_gnt2[6],
    arbout17_gnt2[6], arbout16_gnt2[6], arbout15_gnt2[6], arbout14_gnt2[6],
    arbout13_gnt2[6], arbout12_gnt2[6], arbout11_gnt2[6], arbout10_gnt2[6],
    arbout09_gnt2[6], arbout08_gnt2[6], arbout07_gnt2[6], arbout06_gnt2[6],
    arbout05_gnt2[6], arbout04_gnt2[6], arbout03_gnt2[6], arbout02_gnt2[6],
    arbout01_gnt2[6], arbout00_gnt2[6]};

  assign arbin07_gnt2 = {
    arbout21_gnt2[7], arbout20_gnt2[7], arbout19_gnt2[7], arbout18_gnt2[7],
    arbout17_gnt2[7], arbout16_gnt2[7], arbout15_gnt2[7], arbout14_gnt2[7],
    arbout13_gnt2[7], arbout12_gnt2[7], arbout11_gnt2[7], arbout10_gnt2[7],
    arbout09_gnt2[7], arbout08_gnt2[7], arbout07_gnt2[7], arbout06_gnt2[7],
    arbout05_gnt2[7], arbout04_gnt2[7], arbout03_gnt2[7], arbout02_gnt2[7],
    arbout01_gnt2[7], arbout00_gnt2[7]};

  assign arbin08_gnt2 = {
    arbout21_gnt2[8], arbout20_gnt2[8], arbout19_gnt2[8], arbout18_gnt2[8],
    arbout17_gnt2[8], arbout16_gnt2[8], arbout15_gnt2[8], arbout14_gnt2[8],
    arbout13_gnt2[8], arbout12_gnt2[8], arbout11_gnt2[8], arbout10_gnt2[8],
    arbout09_gnt2[8], arbout08_gnt2[8], arbout07_gnt2[8], arbout06_gnt2[8],
    arbout05_gnt2[8], arbout04_gnt2[8], arbout03_gnt2[8], arbout02_gnt2[8],
    arbout01_gnt2[8], arbout00_gnt2[8]};

  assign arbin09_gnt2 = {
    arbout21_gnt2[9], arbout20_gnt2[9], arbout19_gnt2[9], arbout18_gnt2[9],
    arbout17_gnt2[9], arbout16_gnt2[9], arbout15_gnt2[9], arbout14_gnt2[9],
    arbout13_gnt2[9], arbout12_gnt2[9], arbout11_gnt2[9], arbout10_gnt2[9],
    arbout09_gnt2[9], arbout08_gnt2[9], arbout07_gnt2[9], arbout06_gnt2[9],
    arbout05_gnt2[9], arbout04_gnt2[9], arbout03_gnt2[9], arbout02_gnt2[9],
    arbout01_gnt2[9], arbout00_gnt2[9]};

  assign arbin10_gnt2 = {
    arbout21_gnt2[10], arbout20_gnt2[10], arbout19_gnt2[10], arbout18_gnt2[10],
    arbout17_gnt2[10], arbout16_gnt2[10], arbout15_gnt2[10], arbout14_gnt2[10],
    arbout13_gnt2[10], arbout12_gnt2[10], arbout11_gnt2[10], arbout10_gnt2[10],
    arbout09_gnt2[10], arbout08_gnt2[10], arbout07_gnt2[10], arbout06_gnt2[10],
    arbout05_gnt2[10], arbout04_gnt2[10], arbout03_gnt2[10], arbout02_gnt2[10],
    arbout01_gnt2[10], arbout00_gnt2[10]};

  assign arbin11_gnt2 = {
    arbout21_gnt2[11], arbout20_gnt2[11], arbout19_gnt2[11], arbout18_gnt2[11],
    arbout17_gnt2[11], arbout16_gnt2[11], arbout15_gnt2[11], arbout14_gnt2[11],
    arbout13_gnt2[11], arbout12_gnt2[11], arbout11_gnt2[11], arbout10_gnt2[11],
    arbout09_gnt2[11], arbout08_gnt2[11], arbout07_gnt2[11], arbout06_gnt2[11],
    arbout05_gnt2[11], arbout04_gnt2[11], arbout03_gnt2[11], arbout02_gnt2[11],
    arbout01_gnt2[11], arbout00_gnt2[11]};

  assign arbin12_gnt2 = {
    arbout21_gnt2[12], arbout20_gnt2[12], arbout19_gnt2[12], arbout18_gnt2[12],
    arbout17_gnt2[12], arbout16_gnt2[12], arbout15_gnt2[12], arbout14_gnt2[12],
    arbout13_gnt2[12], arbout12_gnt2[12], arbout11_gnt2[12], arbout10_gnt2[12],
    arbout09_gnt2[12], arbout08_gnt2[12], arbout07_gnt2[12], arbout06_gnt2[12],
    arbout05_gnt2[12], arbout04_gnt2[12], arbout03_gnt2[12], arbout02_gnt2[12],
    arbout01_gnt2[12], arbout00_gnt2[12]};

  assign arbin13_gnt2 = {
    arbout21_gnt2[13], arbout20_gnt2[13], arbout19_gnt2[13], arbout18_gnt2[13],
    arbout17_gnt2[13], arbout16_gnt2[13], arbout15_gnt2[13], arbout14_gnt2[13],
    arbout13_gnt2[13], arbout12_gnt2[13], arbout11_gnt2[13], arbout10_gnt2[13],
    arbout09_gnt2[13], arbout08_gnt2[13], arbout07_gnt2[13], arbout06_gnt2[13],
    arbout05_gnt2[13], arbout04_gnt2[13], arbout03_gnt2[13], arbout02_gnt2[13],
    arbout01_gnt2[13], arbout00_gnt2[13]};

  assign arbin14_gnt2 = {
    arbout21_gnt2[14], arbout20_gnt2[14], arbout19_gnt2[14], arbout18_gnt2[14],
    arbout17_gnt2[14], arbout16_gnt2[14], arbout15_gnt2[14], arbout14_gnt2[14],
    arbout13_gnt2[14], arbout12_gnt2[14], arbout11_gnt2[14], arbout10_gnt2[14],
    arbout09_gnt2[14], arbout08_gnt2[14], arbout07_gnt2[14], arbout06_gnt2[14],
    arbout05_gnt2[14], arbout04_gnt2[14], arbout03_gnt2[14], arbout02_gnt2[14],
    arbout01_gnt2[14], arbout00_gnt2[14]};

  assign arbin15_gnt2 = {
    arbout21_gnt2[15], arbout20_gnt2[15], arbout19_gnt2[15], arbout18_gnt2[15],
    arbout17_gnt2[15], arbout16_gnt2[15], arbout15_gnt2[15], arbout14_gnt2[15],
    arbout13_gnt2[15], arbout12_gnt2[15], arbout11_gnt2[15], arbout10_gnt2[15],
    arbout09_gnt2[15], arbout08_gnt2[15], arbout07_gnt2[15], arbout06_gnt2[15],
    arbout05_gnt2[15], arbout04_gnt2[15], arbout03_gnt2[15], arbout02_gnt2[15],
    arbout01_gnt2[15], arbout00_gnt2[15]};

  assign arbin16_gnt2 = {
    arbout21_gnt2[16], arbout20_gnt2[16], arbout19_gnt2[16], arbout18_gnt2[16],
    arbout17_gnt2[16], arbout16_gnt2[16], arbout15_gnt2[16], arbout14_gnt2[16],
    arbout13_gnt2[16], arbout12_gnt2[16], arbout11_gnt2[16], arbout10_gnt2[16],
    arbout09_gnt2[16], arbout08_gnt2[16], arbout07_gnt2[16], arbout06_gnt2[16],
    arbout05_gnt2[16], arbout04_gnt2[16], arbout03_gnt2[16], arbout02_gnt2[16],
    arbout01_gnt2[16], arbout00_gnt2[16]};

  assign arbin17_gnt2 = {
    arbout21_gnt2[17], arbout20_gnt2[17], arbout19_gnt2[17], arbout18_gnt2[17],
    arbout17_gnt2[17], arbout16_gnt2[17], arbout15_gnt2[17], arbout14_gnt2[17],
    arbout13_gnt2[17], arbout12_gnt2[17], arbout11_gnt2[17], arbout10_gnt2[17],
    arbout09_gnt2[17], arbout08_gnt2[17], arbout07_gnt2[17], arbout06_gnt2[17],
    arbout05_gnt2[17], arbout04_gnt2[17], arbout03_gnt2[17], arbout02_gnt2[17],
    arbout01_gnt2[17], arbout00_gnt2[17]};

  assign arbin18_gnt2 = {
    arbout21_gnt2[18], arbout20_gnt2[18], arbout19_gnt2[18], arbout18_gnt2[18],
    arbout17_gnt2[18], arbout16_gnt2[18], arbout15_gnt2[18], arbout14_gnt2[18],
    arbout13_gnt2[18], arbout12_gnt2[18], arbout11_gnt2[18], arbout10_gnt2[18],
    arbout09_gnt2[18], arbout08_gnt2[18], arbout07_gnt2[18], arbout06_gnt2[18],
    arbout05_gnt2[18], arbout04_gnt2[18], arbout03_gnt2[18], arbout02_gnt2[18],
    arbout01_gnt2[18], arbout00_gnt2[18]};

  assign arbin19_gnt2 = {
    arbout21_gnt2[19], arbout20_gnt2[19], arbout19_gnt2[19], arbout18_gnt2[19],
    arbout17_gnt2[19], arbout16_gnt2[19], arbout15_gnt2[19], arbout14_gnt2[19],
    arbout13_gnt2[19], arbout12_gnt2[19], arbout11_gnt2[19], arbout10_gnt2[19],
    arbout09_gnt2[19], arbout08_gnt2[19], arbout07_gnt2[19], arbout06_gnt2[19],
    arbout05_gnt2[19], arbout04_gnt2[19], arbout03_gnt2[19], arbout02_gnt2[19],
    arbout01_gnt2[19], arbout00_gnt2[19]};

  assign arbin20_gnt2 = {
    arbout21_gnt2[20], arbout20_gnt2[20], arbout19_gnt2[20], arbout18_gnt2[20],
    arbout17_gnt2[20], arbout16_gnt2[20], arbout15_gnt2[20], arbout14_gnt2[20],
    arbout13_gnt2[20], arbout12_gnt2[20], arbout11_gnt2[20], arbout10_gnt2[20],
    arbout09_gnt2[20], arbout08_gnt2[20], arbout07_gnt2[20], arbout06_gnt2[20],
    arbout05_gnt2[20], arbout04_gnt2[20], arbout03_gnt2[20], arbout02_gnt2[20],
    arbout01_gnt2[20], arbout00_gnt2[20]};

  assign arbin21_gnt2 = {
    arbout21_gnt2[21], arbout20_gnt2[21], arbout19_gnt2[21], arbout18_gnt2[21],
    arbout17_gnt2[21], arbout16_gnt2[21], arbout15_gnt2[21], arbout14_gnt2[21],
    arbout13_gnt2[21], arbout12_gnt2[21], arbout11_gnt2[21], arbout10_gnt2[21],
    arbout09_gnt2[21], arbout08_gnt2[21], arbout07_gnt2[21], arbout06_gnt2[21],
    arbout05_gnt2[21], arbout04_gnt2[21], arbout03_gnt2[21], arbout02_gnt2[21],
    arbout01_gnt2[21], arbout00_gnt2[21]};


endmodule
